LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE WORK.ddPackage.ALL;

ENTITY packetParser IS
	PORT (
		clk : IN std_logic;
		packet_in : IN std_logic_vector(7 DOWNTO 0);
		valid_in : IN std_logic:= '0';
		hello_received : OUT std_logic:= '0' ;
		--set i`f hello packet completely received
		dd_received : OUT std_logic:='0';
		-- set if dd packet completely received
		-- respective output ports
		DD : OUT databaseDescription
);
END packetParser;

ARCHITECTURE packetParser_arc OF packetParser IS
--	SIGNAL DD : databaseDescription; 
	SIGNAL counter : std_logic_vector(15 DOWNTO 0) := "0000000000000000";

	SIGNAL version, packetType : std_logic_vector(7 DOWNTO 0):= "00000000";
	SIGNAL packetLength, checksum, auType : std_logic_vector(15 DOWNTO 0);
	SIGNAL routerID, areaID : std_logic_vector(31 DOWNTO 0);
	SIGNAL authentication : std_logic_vector(63 DOWNTO 0);

	SIGNAL networkMask, routerDeadInterval, designatedRouter, backupDesignatedRouter : std_logic_vector(31 DOWNTO 0);
	SIGNAL neighbour1, neighbour2, neighbour3, neighbour4, neighbour5, neighbour6, neighbour7, neighbour8 : std_logic_vector(31 DOWNTO 0);
	SIGNAL helloInterval : std_logic_vector(15 DOWNTO 0);
	SIGNAL options1, rtrPri : std_logic_vector(7 DOWNTO 0);

	SIGNAL zero1, zero2, options2, random : std_logic_vector(7 DOWNTO 0);
	SIGNAL ddSequenceNumber : std_logic_vector(31 DOWNTO 0);
	signal hello_done :std_logic:= '0';

	SIGNAL lsType, linkStateID, advertisingRouter : std_logic_vector(31 DOWNTO 0);

BEGIN
	PROCESS (clk)
	BEGIN
		IF rising_edge(clk) THEN
			IF (valid_in = '1') THEN
				CASE(counter) IS
					WHEN "0000000000000000" =>
					version <= packet_in;
					counter <= "0000000000000001";
					WHEN "0000000000000001" =>
					packetType <= packet_in;
					counter <= "0000000000000010";
					WHEN "0000000000000010" =>
					packetLength(15 DOWNTO 8) <= packet_in;
					counter <= "0000000000000011";
					WHEN "0000000000000011" =>
					packetLength(7 DOWNTO 0) <= packet_in;
					counter <= "0000000000000100";
					WHEN "0000000000000100" =>
					routerID(31 DOWNTO 24) <= packet_in;
					counter <= "0000000000000101";
					WHEN "0000000000000101" =>
					routerID(23 DOWNTO 16) <= packet_in;
					counter <= "0000000000000110";
					WHEN "0000000000000110" =>
					routerID(15 DOWNTO 8) <= packet_in;
					counter <= "0000000000000111";
					WHEN "0000000000000111" =>
					routerID(7 DOWNTO 0) <= packet_in;
					counter <= "0000000000001000";
					WHEN "0000000000001000" =>
					areaID(31 DOWNTO 24) <= packet_in;
					counter <= "0000000000001001";
					WHEN "0000000000001001" =>
					areaID(23 DOWNTO 16) <= packet_in;
					counter <= "0000000000001010";
					WHEN "0000000000001010" =>
					areaID(15 DOWNTO 8) <= packet_in;
					counter <= "0000000000001011";
					WHEN "0000000000001011" =>
					areaID(7 DOWNTO 0) <= packet_in;
					counter <= "0000000000001100";
					WHEN "0000000000001100" =>
					checksum(15 DOWNTO 8) <= packet_in;
					counter <= "0000000000001101";
					WHEN "0000000000001101" =>
					checksum(7 DOWNTO 0) <= packet_in;
					counter <= "0000000000001110";
					WHEN "0000000000001110" =>
					auType(15 DOWNTO 8) <= packet_in;
					counter <= "0000000000001111";
					WHEN "0000000000001111" =>
					auType(7 DOWNTO 0) <= packet_in;
					counter <= "0000000000010000";
					WHEN "0000000000010000" =>
					authentication(63 DOWNTO 56) <= packet_in;
					counter <= "0000000000010001";
					WHEN "0000000000010001" =>
					authentication(55 DOWNTO 48) <= packet_in;
					counter <= "0000000000010010";
					WHEN "0000000000010010" =>
					authentication(47 DOWNTO 40) <= packet_in;
					counter <= "0000000000010011";
					WHEN "0000000000010011" =>
					authentication(39 DOWNTO 32) <= packet_in;
					counter <= "0000000000010100";
					WHEN "0000000000010100" =>
					authentication(31 DOWNTO 24) <= packet_in;
					counter <= "0000000000010101";
					WHEN "0000000000010101" =>
					authentication(23 DOWNTO 16) <= packet_in;
					counter <= "0000000000010110";
					WHEN "0000000000010110" =>
					authentication(15 DOWNTO 8) <= packet_in;
					counter <= "0000000000010111";
					WHEN "0000000000010111" =>
					authentication(7 DOWNTO 0) <= packet_in;
					counter <= "0000000000011000";
					WHEN OTHERS =>
					NULL;
				END CASE;

				CASE(packetType) IS
					when "00000001" =>  -- hello packet begins here
						
						dd_received <= '0';
						case(counter) is
							when "0000000000011000" => 
								networkMask(31 downto 24) <= packet_in;
								counter <= "0000000000011001";
							when "0000000000011001" => 
								networkMask(23 downto 16) <= packet_in;
								counter <= "0000000000011010";
							when "0000000000011010" =>
								networkMask(15 downto 8) <= packet_in; 
								counter <= "0000000000011011";
							when "0000000000011011" => 
								networkMask(7 downto 0) <= packet_in;
								counter <= "0000000000011100";
							when "0000000000011100" => 
								helloInterval(15 downto 8) <= packet_in;
								counter <= "0000000000011101";
							when "0000000000011101" => 
								helloInterval(7 downto 0) <= packet_in;
								counter <= "0000000000011110";
							when "0000000000011110" =>
								options1(7 downto 0) <= packet_in;
								counter <= "0000000000011111";
							when "0000000000011111" =>
								rtrPri(7 downto 0) <= packet_in;
								counter <= "0000000000100000";
							when "0000000000100000" =>
								routerDeadInterval(31 downto 24) <= packet_in;
								counter <= "0000000000100001";
							when "0000000000100001" =>
								routerDeadInterval(23 downto 16) <= packet_in;
								counter <= "0000000000100010";
							when "0000000000100010" =>
								routerDeadInterval(15 downto 8) <= packet_in;
								counter <= "0000000000100011";
							when "0000000000100011" =>
								routerDeadInterval(7 downto 0) <= packet_in;
								counter <= "0000000000100100";
							when "0000000000100100" =>
								designatedRouter(31 downto 24) <= packet_in;
								counter <= "0000000000100101";
							when "0000000000100101" =>
								designatedRouter(23 downto 16) <= packet_in;
								counter <= "0000000000100110";
							when "0000000000100110" =>
								designatedRouter(15 downto 8) <= packet_in;
								counter <= "0000000000100111";
							when "0000000000100111" =>
								designatedRouter(7 downto 0) <= packet_in;
								counter <= "0000000000101000";
							when "0000000000101000" =>
								backupDesignatedRouter(31 downto 24) <= packet_in;
								counter <= "0000000000101001";
							when "0000000000101001" =>
								backupDesignatedRouter(23 downto 16) <= packet_in;
								counter <= "0000000000101010";
							when "0000000000101010" =>
								backupDesignatedRouter(15 downto 8) <= packet_in;
								counter <= "0000000000101011";
							when "0000000000101011" =>
								backupDesignatedRouter(7 downto 0) <= packet_in;
								counter <= "0000000000101100";

									 when "0000000000101100" =>
                                neighbour1(31 downto 24) <= packet_in;
                                counter <= "0000000000101101";
                            when "0000000000101101" =>
                                neighbour1(23 downto 16) <= packet_in;
                                counter <= "0000000000101110";
                            when "0000000000101110" =>
                                neighbour1(15 downto 8) <= packet_in;
                                counter <= "0000000000101111";
                            when "0000000000101111" =>
                                neighbour1(7 downto 0) <= packet_in;
                                counter <= "0000000000110000";
                            when "0000000000110000" =>
                                neighbour2(31 downto 24) <= packet_in;
                                counter <= "0000000000110001";
                            when "0000000000110001" =>
                                neighbour2(23 downto 16) <= packet_in;
                                counter <= "0000000000110010";
                            when "0000000000110010" =>
                                neighbour2(15 downto 8) <= packet_in;
                                counter <= "0000000000110011";
                            when "0000000000110011" =>
                                neighbour2(7 downto 0) <= packet_in;
                                counter <= "0000000000110100";
                            when "0000000000110100" =>
                                neighbour3(31 downto 24) <= packet_in;
                                counter <= "0000000000110101";
                            when "0000000000110101" =>
                                neighbour3(23 downto 16) <= packet_in;
                                counter <= "0000000000110110";
                            when "0000000000110110" =>
                                neighbour3(15 downto 8) <= packet_in;
                                counter <= "0000000000110111";
                            when "0000000000110111" =>
                                neighbour3(7 downto 0) <= packet_in;
                                counter <= "0000000000111000";
                            when "0000000000111000" =>
                                neighbour4(31 downto 24) <= packet_in;
                                counter <= "0000000000111001";
                            when "0000000000111001" =>
                                neighbour4(23 downto 16) <= packet_in;
                                counter <= "0000000000111010";
                            when "0000000000111010" =>
                                neighbour4(15 downto 8) <= packet_in;
                                counter <= "0000000000111011";
                            when "0000000000111011" =>
                                neighbour4(7 downto 0) <= packet_in;
                                counter <= "0000000000111100";
                            when "0000000000111100" =>
                                neighbour5(31 downto 24) <= packet_in;
                                counter <= "0000000000111101";
                            when "0000000000111101" =>
                                neighbour5(23 downto 16) <= packet_in;
                                counter <= "0000000000111110";
                            when "0000000000111110" =>
                                neighbour5(15 downto 8) <= packet_in;
                                counter <= "0000000000111111";
                            when "0000000000111111" =>
                                neighbour5(7 downto 0) <= packet_in;
                                counter <= "0000000001000000";
                            when "0000000001000000" =>
                                neighbour6(31 downto 24) <= packet_in;
                                counter <= "0000000001000001";
                            when "0000000001000001" =>
                                neighbour6(23 downto 16) <= packet_in;
                                counter <= "0000000001000010";
                            when "0000000001000010" =>
                                neighbour6(15 downto 8) <= packet_in;
                                counter <= "0000000001000011";
                            when "0000000001000011" =>
                                neighbour6(7 downto 0) <= packet_in;
                                counter <= "0000000001000100";
                            when "0000000001000100" =>
                                neighbour7(31 downto 24) <= packet_in;
                                counter <= "0000000001000101";
                            when "0000000001000101" =>
                                neighbour7(23 downto 16) <= packet_in;
                                counter <= "0000000001000110";
                            when "0000000001000110" =>
                                neighbour7(15 downto 8) <= packet_in;
                                counter <= "0000000001000111";
                            when "0000000001000111" =>
                                neighbour7(7 downto 0) <= packet_in;
                                counter <= "0000000001001000";
                            when "0000000001001000" =>
                                neighbour8(31 downto 24) <= packet_in;
                                counter <= "0000000001001001";
                            when "0000000001001001" =>
                                neighbour8(23 downto 16) <= packet_in;
                                counter <= "0000000001001010";
                            when "0000000001001010" =>
                                neighbour8(15 downto 8) <= packet_in;
                                counter <= "0000000001001011";
                            when "0000000001001011" =>
                                neighbour8(7 downto 0) <= packet_in;
										  hello_received <= '1';        
										counter <= "0000000000000000";
--											hello_done <= '1';
--									 when "0000000001001100" =>
--									 	  report "Hail satan";
--										  hello_received <= '1';        
--										  counter <= "0000000000000000";
                            when others =>
                                null;
								end case; -- case for hello packet ends here
					WHEN "00000010" => 					-- case for database description packet begins here
						hello_received <= '0';
					  report "Hail satan 2";

					CASE(counter) IS
						WHEN "0000000000011000" =>
						zero1(7 DOWNTO 0) <= packet_in;
						counter <= "0000000000011001";
						WHEN "0000000000011001" =>
						zero2(7 DOWNTO 0) <= packet_in;
						counter <= "0000000000011010";
						WHEN "0000000000011010" =>
						options2(7 DOWNTO 0) <= packet_in;
						counter <= "0000000000011011";
						WHEN "0000000000011011" =>
						random(7 DOWNTO 0) <= packet_in;
						counter <= "0000000000011100";
						WHEN "0000000000011100" =>
						ddSequenceNumber(31 DOWNTO 24) <= packet_in;
						counter <= "0000000000011101";
						WHEN "0000000000011101" =>
						ddSequenceNumber(23 DOWNTO 16) <= packet_in;
						counter <= "0000000000011110";
						WHEN "0000000000011110" =>
						ddSequenceNumber(15 DOWNTO 8) <= packet_in;
						counter <= "0000000000011111";
						WHEN "0000000000011111" =>
						ddSequenceNumber(7 DOWNTO 0) <= packet_in;
						counter <= "0000000000100000";
						-- till here, the whole packet is parsed according to the standard,
						-- now the 32 link state advertisements will be read and stored in 
						-- an array of size 32 X 92 , where 92 is the size of one advertisement
						WHEN "0000000000100000" =>
						DD(0,0) <= packet_in;
						counter <= "0000000000100001";
						WHEN "0000000000100001" =>
						DD(0,1) <= packet_in;
						counter <= "0000000000100010";
						WHEN "0000000000100010" =>
						DD(0,2) <= packet_in;
						counter <= "0000000000100011";
						WHEN "0000000000100011" =>
						DD(0,3) <= packet_in;
						counter <= "0000000000100100";
						WHEN "0000000000100100" =>
						DD(0,4) <= packet_in;
						counter <= "0000000000100101";
						WHEN "0000000000100101" =>
						DD(0, 5) <= packet_in;
						counter <= "0000000000100110";
						WHEN "0000000000100110" =>
						DD(0, 6) <= packet_in;
						counter <= "0000000000100111";
						WHEN "0000000000100111" =>
						DD(0, 7) <= packet_in;
						counter <= "0000000000101000";
						WHEN "0000000000101000" =>
						DD(0, 8) <= packet_in;
						counter <= "0000000000101001";
						WHEN "0000000000101001" =>
						DD(0, 9) <= packet_in;
						counter <= "0000000000101010";
						WHEN "0000000000101010" =>
						DD(0, 10) <= packet_in;
						counter <= "0000000000101011";
						WHEN "0000000000101011" =>
						DD(0, 11) <= packet_in;
						counter <= "0000000000101100";
						WHEN "0000000000101100" =>
						DD(0, 12) <= packet_in;
						counter <= "0000000000101101";
						WHEN "0000000000101101" =>
						DD(0, 13) <= packet_in;
						counter <= "0000000000101110";
						WHEN "0000000000101110" =>
						DD(0, 14) <= packet_in;
						counter <= "0000000000101111";
						WHEN "0000000000101111" =>
						DD(0, 15) <= packet_in;
						counter <= "0000000000110000";
						WHEN "0000000000110000" =>
						DD(0, 16) <= packet_in;
						counter <= "0000000000110001";
						WHEN "0000000000110001" =>
						DD(0, 17) <= packet_in;
						counter <= "0000000000110010";
						WHEN "0000000000110010" =>
						DD(0, 18) <= packet_in;
						counter <= "0000000000110011";
						WHEN "0000000000110011" =>
						DD(0, 19) <= packet_in;
						counter <= "0000000000110100";
						WHEN "0000000000110100" =>
						DD(0, 20) <= packet_in;
						counter <= "0000000000110101";
						WHEN "0000000000110101" =>
						DD(0, 21) <= packet_in;
						counter <= "0000000000110110";
						WHEN "0000000000110110" =>
						DD(0, 22) <= packet_in;
						counter <= "0000000000110111";
						WHEN "0000000000110111" =>
						DD(0, 23) <= packet_in;
						counter <= "0000000000111000";
						WHEN "0000000000111000" =>
						DD(0, 24) <= packet_in;
						counter <= "0000000000111001";
						WHEN "0000000000111001" =>
						DD(0, 25) <= packet_in;
						counter <= "0000000000111010";
						WHEN "0000000000111010" =>
						DD(0, 26) <= packet_in;
						counter <= "0000000000111011";
						WHEN "0000000000111011" =>
						DD(0, 27) <= packet_in;
						counter <= "0000000000111100";
						WHEN "0000000000111100" =>
						DD(0, 28) <= packet_in;
						counter <= "0000000000111101";
						WHEN "0000000000111101" =>
						DD(0, 29) <= packet_in;
						counter <= "0000000000111110";
						WHEN "0000000000111110" =>
						DD(0, 30) <= packet_in;
						counter <= "0000000000111111";
						WHEN "0000000000111111" =>
						DD(0, 31) <= packet_in;
						counter <= "0000000001000000";
						WHEN "0000000001000000" =>
						DD(0, 32) <= packet_in;
						counter <= "0000000001000001";
						WHEN "0000000001000001" =>
						DD(0, 33) <= packet_in;
						counter <= "0000000001000010";
						WHEN "0000000001000010" =>
						DD(0, 34) <= packet_in;
						counter <= "0000000001000011";
						WHEN "0000000001000011" =>
						DD(0, 35) <= packet_in;
						counter <= "0000000001000100";
						WHEN "0000000001000100" =>
						DD(0, 36) <= packet_in;
						counter <= "0000000001000101";
						WHEN "0000000001000101" =>
						DD(0, 37) <= packet_in;
						counter <= "0000000001000110";
						WHEN "0000000001000110" =>
						DD(0, 38) <= packet_in;
						counter <= "0000000001000111";
						WHEN "0000000001000111" =>
						DD(0, 39) <= packet_in;
						counter <= "0000000001001000";
						WHEN "0000000001001000" =>
						DD(0, 40) <= packet_in;
						counter <= "0000000001001001";
						WHEN "0000000001001001" =>
						DD(0, 41) <= packet_in;
						counter <= "0000000001001010";
						WHEN "0000000001001010" =>
						DD(0, 42) <= packet_in;
						counter <= "0000000001001011";
						WHEN "0000000001001011" =>
						DD(0, 43) <= packet_in;
						counter <= "0000000001001100";
						WHEN "0000000001001100" =>
						DD(0, 44) <= packet_in;
						counter <= "0000000001001101";
						WHEN "0000000001001101" =>
						DD(0, 45) <= packet_in;
						counter <= "0000000001001110";
						WHEN "0000000001001110" =>
						DD(0, 46) <= packet_in;
						counter <= "0000000001001111";
						WHEN "0000000001001111" =>
						DD(0, 47) <= packet_in;
						counter <= "0000000001010000";
						WHEN "0000000001010000" =>
						DD(0, 48) <= packet_in;
						counter <= "0000000001010001";
						WHEN "0000000001010001" =>
						DD(0, 49) <= packet_in;
						counter <= "0000000001010010";
						WHEN "0000000001010010" =>
						DD(0, 50) <= packet_in;
						counter <= "0000000001010011";
						WHEN "0000000001010011" =>
						DD(0, 51) <= packet_in;
						counter <= "0000000001010100";
						WHEN "0000000001010100" =>
						DD(0, 52) <= packet_in;
						counter <= "0000000001010101";
						WHEN "0000000001010101" =>
						DD(0, 53) <= packet_in;
						counter <= "0000000001010110";
						WHEN "0000000001010110" =>
						DD(0, 54) <= packet_in;
						counter <= "0000000001010111";
						WHEN "0000000001010111" =>
						DD(0, 55) <= packet_in;
						counter <= "0000000001011000";
						WHEN "0000000001011000" =>
						DD(0, 56) <= packet_in;
						counter <= "0000000001011001";
						WHEN "0000000001011001" =>
						DD(0, 57) <= packet_in;
						counter <= "0000000001011010";
						WHEN "0000000001011010" =>
						DD(0, 58) <= packet_in;
						counter <= "0000000001011011";
						WHEN "0000000001011011" =>
						DD(0, 59) <= packet_in;
						counter <= "0000000001011100";
						WHEN "0000000001011100" =>
						DD(0, 60) <= packet_in;
						counter <= "0000000001011101";
						WHEN "0000000001011101" =>
						DD(0, 61) <= packet_in;
						counter <= "0000000001011110";
						WHEN "0000000001011110" =>
						DD(0, 62) <= packet_in;
						counter <= "0000000001011111";
						WHEN "0000000001011111" =>
						DD(0, 63) <= packet_in;
						counter <= "0000000001100000";
						WHEN "0000000001100000" =>
						DD(0, 64) <= packet_in;
						counter <= "0000000001100001";
						WHEN "0000000001100001" =>
						DD(0, 65) <= packet_in;
						counter <= "0000000001100010";
						WHEN "0000000001100010" =>
						DD(0, 66) <= packet_in;
						counter <= "0000000001100011";
						WHEN "0000000001100011" =>
						DD(0, 67) <= packet_in;
						counter <= "0000000001100100";
						WHEN "0000000001100100" =>
						DD(0, 68) <= packet_in;
						counter <= "0000000001100101";
						WHEN "0000000001100101" =>
						DD(0, 69) <= packet_in;
						counter <= "0000000001100110";
						WHEN "0000000001100110" =>
						DD(0, 70) <= packet_in;
						counter <= "0000000001100111";
						WHEN "0000000001100111" =>
						DD(0, 71) <= packet_in;
						counter <= "0000000001101000";
						WHEN "0000000001101000" =>
						DD(0, 72) <= packet_in;
						counter <= "0000000001101001";
						WHEN "0000000001101001" =>
						DD(0, 73) <= packet_in;
						counter <= "0000000001101010";
						WHEN "0000000001101010" =>
						DD(0, 74) <= packet_in;
						counter <= "0000000001101011";
						WHEN "0000000001101011" =>
						DD(0, 75) <= packet_in;
						counter <= "0000000001101100";
						WHEN "0000000001101100" =>
						DD(0, 76) <= packet_in;
						counter <= "0000000001101101";
						WHEN "0000000001101101" =>
						DD(0, 77) <= packet_in;
						counter <= "0000000001101110";
						WHEN "0000000001101110" =>
						DD(0, 78) <= packet_in;
						counter <= "0000000001101111";
						WHEN "0000000001101111" =>
						DD(0, 79) <= packet_in;
						counter <= "0000000001110000";
						WHEN "0000000001110000" =>
						DD(0, 80) <= packet_in;
						counter <= "0000000001110001";
						WHEN "0000000001110001" =>
						DD(0, 81) <= packet_in;
						counter <= "0000000001110010";
						WHEN "0000000001110010" =>
						DD(0, 82) <= packet_in;
						counter <= "0000000001110011";
						WHEN "0000000001110011" =>
						DD(0, 83) <= packet_in;
						counter <= "0000000001110100";
						WHEN "0000000001110100" =>
						DD(0, 84) <= packet_in;
						counter <= "0000000001110101";
						WHEN "0000000001110101" =>
						DD(0, 85) <= packet_in;
						counter <= "0000000001110110";
						WHEN "0000000001110110" =>
						DD(0, 86) <= packet_in;
						counter <= "0000000001110111";
						WHEN "0000000001110111" =>
						DD(0, 87) <= packet_in;
						counter <= "0000000001111000";
						WHEN "0000000001111000" =>
						DD(0, 88) <= packet_in;
						counter <= "0000000001111001";
						WHEN "0000000001111001" =>
						DD(0, 89) <= packet_in;
						counter <= "0000000001111010";
						WHEN "0000000001111010" =>
						DD(0, 90) <= packet_in;
						counter <= "0000000001111011";
						WHEN "0000000001111011" =>
						DD(0, 91) <= packet_in;
						counter <= "0000000001111100";
						WHEN "0000000001111100" =>
						DD(1, 0) <= packet_in;
						counter <= "0000000001111101";
						WHEN "0000000001111101" =>
						DD(1, 1) <= packet_in;
						counter <= "0000000001111110";
						WHEN "0000000001111110" =>
						DD(1, 2) <= packet_in;
						counter <= "0000000001111111";
						WHEN "0000000001111111" =>
						DD(1, 3) <= packet_in;
						counter <= "0000000010000000";
						WHEN "0000000010000000" =>
						DD(1, 4) <= packet_in;
						counter <= "0000000010000001";
						WHEN "0000000010000001" =>
						DD(1, 5) <= packet_in;
						counter <= "0000000010000010";
						WHEN "0000000010000010" =>
						DD(1, 6) <= packet_in;
						counter <= "0000000010000011";
						WHEN "0000000010000011" =>
						DD(1, 7) <= packet_in;
						counter <= "0000000010000100";
						WHEN "0000000010000100" =>
						DD(1, 8) <= packet_in;
						counter <= "0000000010000101";
						WHEN "0000000010000101" =>
						DD(1, 9) <= packet_in;
						counter <= "0000000010000110";
						WHEN "0000000010000110" =>
						DD(1, 10) <= packet_in;
						counter <= "0000000010000111";
						WHEN "0000000010000111" =>
						DD(1, 11) <= packet_in;
						counter <= "0000000010001000";
						WHEN "0000000010001000" =>
						DD(1, 12) <= packet_in;
						counter <= "0000000010001001";
						WHEN "0000000010001001" =>
						DD(1, 13) <= packet_in;
						counter <= "0000000010001010";
						WHEN "0000000010001010" =>
						DD(1, 14) <= packet_in;
						counter <= "0000000010001011";
						WHEN "0000000010001011" =>
						DD(1, 15) <= packet_in;
						counter <= "0000000010001100";
						WHEN "0000000010001100" =>
						DD(1, 16) <= packet_in;
						counter <= "0000000010001101";
						WHEN "0000000010001101" =>
						DD(1, 17) <= packet_in;
						counter <= "0000000010001110";
						WHEN "0000000010001110" =>
						DD(1, 18) <= packet_in;
						counter <= "0000000010001111";
						WHEN "0000000010001111" =>
						DD(1, 19) <= packet_in;
						counter <= "0000000010010000";
						WHEN "0000000010010000" =>
						DD(1, 20) <= packet_in;
						counter <= "0000000010010001";
						WHEN "0000000010010001" =>
						DD(1, 21) <= packet_in;
						counter <= "0000000010010010";
						WHEN "0000000010010010" =>
						DD(1, 22) <= packet_in;
						counter <= "0000000010010011";
						WHEN "0000000010010011" =>
						DD(1, 23) <= packet_in;
						counter <= "0000000010010100";
						WHEN "0000000010010100" =>
						DD(1, 24) <= packet_in;
						counter <= "0000000010010101";
						WHEN "0000000010010101" =>
						DD(1, 25) <= packet_in;
						counter <= "0000000010010110";
						WHEN "0000000010010110" =>
						DD(1, 26) <= packet_in;
						counter <= "0000000010010111";
						WHEN "0000000010010111" =>
						DD(1, 27) <= packet_in;
						counter <= "0000000010011000";
						WHEN "0000000010011000" =>
						DD(1, 28) <= packet_in;
						counter <= "0000000010011001";
						WHEN "0000000010011001" =>
						DD(1, 29) <= packet_in;
						counter <= "0000000010011010";
						WHEN "0000000010011010" =>
						DD(1, 30) <= packet_in;
						counter <= "0000000010011011";
						WHEN "0000000010011011" =>
						DD(1, 31) <= packet_in;
						counter <= "0000000010011100";
						WHEN "0000000010011100" =>
						DD(1, 32) <= packet_in;
						counter <= "0000000010011101";
						WHEN "0000000010011101" =>
						DD(1, 33) <= packet_in;
						counter <= "0000000010011110";
						WHEN "0000000010011110" =>
						DD(1, 34) <= packet_in;
						counter <= "0000000010011111";
						WHEN "0000000010011111" =>
						DD(1, 35) <= packet_in;
						counter <= "0000000010100000";
						WHEN "0000000010100000" =>
						DD(1, 36) <= packet_in;
						counter <= "0000000010100001";
						WHEN "0000000010100001" =>
						DD(1, 37) <= packet_in;
						counter <= "0000000010100010";
						WHEN "0000000010100010" =>
						DD(1, 38) <= packet_in;
						counter <= "0000000010100011";
						WHEN "0000000010100011" =>
						DD(1, 39) <= packet_in;
						counter <= "0000000010100100";
						WHEN "0000000010100100" =>
						DD(1, 40) <= packet_in;
						counter <= "0000000010100101";
						WHEN "0000000010100101" =>
						DD(1, 41) <= packet_in;
						counter <= "0000000010100110";
						WHEN "0000000010100110" =>
						DD(1, 42) <= packet_in;
						counter <= "0000000010100111";
						WHEN "0000000010100111" =>
						DD(1, 43) <= packet_in;
						counter <= "0000000010101000";
						WHEN "0000000010101000" =>
						DD(1, 44) <= packet_in;
						counter <= "0000000010101001";
						WHEN "0000000010101001" =>
						DD(1, 45) <= packet_in;
						counter <= "0000000010101010";
						WHEN "0000000010101010" =>
						DD(1, 46) <= packet_in;
						counter <= "0000000010101011";
						WHEN "0000000010101011" =>
						DD(1, 47) <= packet_in;
						counter <= "0000000010101100";
						WHEN "0000000010101100" =>
						DD(1, 48) <= packet_in;
						counter <= "0000000010101101";
						WHEN "0000000010101101" =>
						DD(1, 49) <= packet_in;
						counter <= "0000000010101110";
						WHEN "0000000010101110" =>
						DD(1, 50) <= packet_in;
						counter <= "0000000010101111";
						WHEN "0000000010101111" =>
						DD(1, 51) <= packet_in;
						counter <= "0000000010110000";
						WHEN "0000000010110000" =>
						DD(1, 52) <= packet_in;
						counter <= "0000000010110001";
						WHEN "0000000010110001" =>
						DD(1, 53) <= packet_in;
						counter <= "0000000010110010";
						WHEN "0000000010110010" =>
						DD(1, 54) <= packet_in;
						counter <= "0000000010110011";
						WHEN "0000000010110011" =>
						DD(1, 55) <= packet_in;
						counter <= "0000000010110100";
						WHEN "0000000010110100" =>
						DD(1, 56) <= packet_in;
						counter <= "0000000010110101";
						WHEN "0000000010110101" =>
						DD(1, 57) <= packet_in;
						counter <= "0000000010110110";
						WHEN "0000000010110110" =>
						DD(1, 58) <= packet_in;
						counter <= "0000000010110111";
						WHEN "0000000010110111" =>
						DD(1, 59) <= packet_in;
						counter <= "0000000010111000";
						WHEN "0000000010111000" =>
						DD(1, 60) <= packet_in;
						counter <= "0000000010111001";
						WHEN "0000000010111001" =>
						DD(1, 61) <= packet_in;
						counter <= "0000000010111010";
						WHEN "0000000010111010" =>
						DD(1, 62) <= packet_in;
						counter <= "0000000010111011";
						WHEN "0000000010111011" =>
						DD(1, 63) <= packet_in;
						counter <= "0000000010111100";
						WHEN "0000000010111100" =>
						DD(1, 64) <= packet_in;
						counter <= "0000000010111101";
						WHEN "0000000010111101" =>
						DD(1, 65) <= packet_in;
						counter <= "0000000010111110";
						WHEN "0000000010111110" =>
						DD(1, 66) <= packet_in;
						counter <= "0000000010111111";
						WHEN "0000000010111111" =>
						DD(1, 67) <= packet_in;
						counter <= "0000000011000000";
						WHEN "0000000011000000" =>
						DD(1, 68) <= packet_in;
						counter <= "0000000011000001";
						WHEN "0000000011000001" =>
						DD(1, 69) <= packet_in;
						counter <= "0000000011000010";
						WHEN "0000000011000010" =>
						DD(1, 70) <= packet_in;
						counter <= "0000000011000011";
						WHEN "0000000011000011" =>
						DD(1, 71) <= packet_in;
						counter <= "0000000011000100";
						WHEN "0000000011000100" =>
						DD(1, 72) <= packet_in;
						counter <= "0000000011000101";
						WHEN "0000000011000101" =>
						DD(1, 73) <= packet_in;
						counter <= "0000000011000110";
						WHEN "0000000011000110" =>
						DD(1, 74) <= packet_in;
						counter <= "0000000011000111";
						WHEN "0000000011000111" =>
						DD(1, 75) <= packet_in;
						counter <= "0000000011001000";
						WHEN "0000000011001000" =>
						DD(1, 76) <= packet_in;
						counter <= "0000000011001001";
						WHEN "0000000011001001" =>
						DD(1, 77) <= packet_in;
						counter <= "0000000011001010";
						WHEN "0000000011001010" =>
						DD(1, 78) <= packet_in;
						counter <= "0000000011001011";
						WHEN "0000000011001011" =>
						DD(1, 79) <= packet_in;
						counter <= "0000000011001100";
						WHEN "0000000011001100" =>
						DD(1, 80) <= packet_in;
						counter <= "0000000011001101";
						WHEN "0000000011001101" =>
						DD(1, 81) <= packet_in;
						counter <= "0000000011001110";
						WHEN "0000000011001110" =>
						DD(1, 82) <= packet_in;
						counter <= "0000000011001111";
						WHEN "0000000011001111" =>
						DD(1, 83) <= packet_in;
						counter <= "0000000011010000";
						WHEN "0000000011010000" =>
						DD(1, 84) <= packet_in;
						counter <= "0000000011010001";
						WHEN "0000000011010001" =>
						DD(1, 85) <= packet_in;
						counter <= "0000000011010010";
						WHEN "0000000011010010" =>
						DD(1, 86) <= packet_in;
						counter <= "0000000011010011";
						WHEN "0000000011010011" =>
						DD(1, 87) <= packet_in;
						counter <= "0000000011010100";
						WHEN "0000000011010100" =>
						DD(1, 88) <= packet_in;
						counter <= "0000000011010101";
						WHEN "0000000011010101" =>
						DD(1, 89) <= packet_in;
						counter <= "0000000011010110";
						WHEN "0000000011010110" =>
						DD(1, 90) <= packet_in;
						counter <= "0000000011010111";
						WHEN "0000000011010111" =>
						DD(1, 91) <= packet_in;
						counter <= "0000000011011000";
						WHEN "0000000011011000" =>
						DD(2, 0) <= packet_in;
						counter <= "0000000011011001";
						WHEN "0000000011011001" =>
						DD(2, 1) <= packet_in;
						counter <= "0000000011011010";
						WHEN "0000000011011010" =>
						DD(2, 2) <= packet_in;
						counter <= "0000000011011011";
						WHEN "0000000011011011" =>
						DD(2, 3) <= packet_in;
						counter <= "0000000011011100";
						WHEN "0000000011011100" =>
						DD(2, 4) <= packet_in;
						counter <= "0000000011011101";
						WHEN "0000000011011101" =>
						DD(2, 5) <= packet_in;
						counter <= "0000000011011110";
						WHEN "0000000011011110" =>
						DD(2, 6) <= packet_in;
						counter <= "0000000011011111";
						WHEN "0000000011011111" =>
						DD(2, 7) <= packet_in;
						counter <= "0000000011100000";
						WHEN "0000000011100000" =>
						DD(2, 8) <= packet_in;
						counter <= "0000000011100001";
						WHEN "0000000011100001" =>
						DD(2, 9) <= packet_in;
						counter <= "0000000011100010";
						WHEN "0000000011100010" =>
						DD(2, 10) <= packet_in;
						counter <= "0000000011100011";
						WHEN "0000000011100011" =>
						DD(2, 11) <= packet_in;
						counter <= "0000000011100100";
						WHEN "0000000011100100" =>
						DD(2, 12) <= packet_in;
						counter <= "0000000011100101";
						WHEN "0000000011100101" =>
						DD(2, 13) <= packet_in;
						counter <= "0000000011100110";
						WHEN "0000000011100110" =>
						DD(2, 14) <= packet_in;
						counter <= "0000000011100111";
						WHEN "0000000011100111" =>
						DD(2, 15) <= packet_in;
						counter <= "0000000011101000";
						WHEN "0000000011101000" =>
						DD(2, 16) <= packet_in;
						counter <= "0000000011101001";
						WHEN "0000000011101001" =>
						DD(2, 17) <= packet_in;
						counter <= "0000000011101010";
						WHEN "0000000011101010" =>
						DD(2, 18) <= packet_in;
						counter <= "0000000011101011";
						WHEN "0000000011101011" =>
						DD(2, 19) <= packet_in;
						counter <= "0000000011101100";
						WHEN "0000000011101100" =>
						DD(2, 20) <= packet_in;
						counter <= "0000000011101101";
						WHEN "0000000011101101" =>
						DD(2, 21) <= packet_in;
						counter <= "0000000011101110";
						WHEN "0000000011101110" =>
						DD(2, 22) <= packet_in;
						counter <= "0000000011101111";
						WHEN "0000000011101111" =>
						DD(2, 23) <= packet_in;
						counter <= "0000000011110000";
						WHEN "0000000011110000" =>
						DD(2, 24) <= packet_in;
						counter <= "0000000011110001";
						WHEN "0000000011110001" =>
						DD(2, 25) <= packet_in;
						counter <= "0000000011110010";
						WHEN "0000000011110010" =>
						DD(2, 26) <= packet_in;
						counter <= "0000000011110011";
						WHEN "0000000011110011" =>
						DD(2, 27) <= packet_in;
						counter <= "0000000011110100";
						WHEN "0000000011110100" =>
						DD(2, 28) <= packet_in;
						counter <= "0000000011110101";
						WHEN "0000000011110101" =>
						DD(2, 29) <= packet_in;
						counter <= "0000000011110110";
						WHEN "0000000011110110" =>
						DD(2, 30) <= packet_in;
						counter <= "0000000011110111";
						WHEN "0000000011110111" =>
						DD(2, 31) <= packet_in;
						counter <= "0000000011111000";
						WHEN "0000000011111000" =>
						DD(2, 32) <= packet_in;
						counter <= "0000000011111001";
						WHEN "0000000011111001" =>
						DD(2, 33) <= packet_in;
						counter <= "0000000011111010";
						WHEN "0000000011111010" =>
						DD(2, 34) <= packet_in;
						counter <= "0000000011111011";
						WHEN "0000000011111011" =>
						DD(2, 35) <= packet_in;
						counter <= "0000000011111100";
						WHEN "0000000011111100" =>
						DD(2, 36) <= packet_in;
						counter <= "0000000011111101";
						WHEN "0000000011111101" =>
						DD(2, 37) <= packet_in;
						counter <= "0000000011111110";
						WHEN "0000000011111110" =>
						DD(2, 38) <= packet_in;
						counter <= "0000000011111111";
						WHEN "0000000011111111" =>
						DD(2, 39) <= packet_in;
						counter <= "0000000100000000";
						WHEN "0000000100000000" =>
						DD(2, 40) <= packet_in;
						counter <= "0000000100000001";
						WHEN "0000000100000001" =>
						DD(2, 41) <= packet_in;
						counter <= "0000000100000010";
						WHEN "0000000100000010" =>
						DD(2, 42) <= packet_in;
						counter <= "0000000100000011";
						WHEN "0000000100000011" =>
						DD(2, 43) <= packet_in;
						counter <= "0000000100000100";
						WHEN "0000000100000100" =>
						DD(2, 44) <= packet_in;
						counter <= "0000000100000101";
						WHEN "0000000100000101" =>
						DD(2, 45) <= packet_in;
						counter <= "0000000100000110";
						WHEN "0000000100000110" =>
						DD(2, 46) <= packet_in;
						counter <= "0000000100000111";
						WHEN "0000000100000111" =>
						DD(2, 47) <= packet_in;
						counter <= "0000000100001000";
						WHEN "0000000100001000" =>
						DD(2, 48) <= packet_in;
						counter <= "0000000100001001";
						WHEN "0000000100001001" =>
						DD(2, 49) <= packet_in;
						counter <= "0000000100001010";
						WHEN "0000000100001010" =>
						DD(2, 50) <= packet_in;
						counter <= "0000000100001011";
						WHEN "0000000100001011" =>
						DD(2, 51) <= packet_in;
						counter <= "0000000100001100";
						WHEN "0000000100001100" =>
						DD(2, 52) <= packet_in;
						counter <= "0000000100001101";
						WHEN "0000000100001101" =>
						DD(2, 53) <= packet_in;
						counter <= "0000000100001110";
						WHEN "0000000100001110" =>
						DD(2, 54) <= packet_in;
						counter <= "0000000100001111";
						WHEN "0000000100001111" =>
						DD(2, 55) <= packet_in;
						counter <= "0000000100010000";
						WHEN "0000000100010000" =>
						DD(2, 56) <= packet_in;
						counter <= "0000000100010001";
						WHEN "0000000100010001" =>
						DD(2, 57) <= packet_in;
						counter <= "0000000100010010";
						WHEN "0000000100010010" =>
						DD(2, 58) <= packet_in;
						counter <= "0000000100010011";
						WHEN "0000000100010011" =>
						DD(2, 59) <= packet_in;
						counter <= "0000000100010100";
						WHEN "0000000100010100" =>
						DD(2, 60) <= packet_in;
						counter <= "0000000100010101";
						WHEN "0000000100010101" =>
						DD(2, 61) <= packet_in;
						counter <= "0000000100010110";
						WHEN "0000000100010110" =>
						DD(2, 62) <= packet_in;
						counter <= "0000000100010111";
						WHEN "0000000100010111" =>
						DD(2, 63) <= packet_in;
						counter <= "0000000100011000";
						WHEN "0000000100011000" =>
						DD(2, 64) <= packet_in;
						counter <= "0000000100011001";
						WHEN "0000000100011001" =>
						DD(2, 65) <= packet_in;
						counter <= "0000000100011010";
						WHEN "0000000100011010" =>
						DD(2, 66) <= packet_in;
						counter <= "0000000100011011";
						WHEN "0000000100011011" =>
						DD(2, 67) <= packet_in;
						counter <= "0000000100011100";
						WHEN "0000000100011100" =>
						DD(2, 68) <= packet_in;
						counter <= "0000000100011101";
						WHEN "0000000100011101" =>
						DD(2, 69) <= packet_in;
						counter <= "0000000100011110";
						WHEN "0000000100011110" =>
						DD(2, 70) <= packet_in;
						counter <= "0000000100011111";
						WHEN "0000000100011111" =>
						DD(2, 71) <= packet_in;
						counter <= "0000000100100000";
						WHEN "0000000100100000" =>
						DD(2, 72) <= packet_in;
						counter <= "0000000100100001";
						WHEN "0000000100100001" =>
						DD(2, 73) <= packet_in;
						counter <= "0000000100100010";
						WHEN "0000000100100010" =>
						DD(2, 74) <= packet_in;
						counter <= "0000000100100011";
						WHEN "0000000100100011" =>
						DD(2, 75) <= packet_in;
						counter <= "0000000100100100";
						WHEN "0000000100100100" =>
						DD(2, 76) <= packet_in;
						counter <= "0000000100100101";
						WHEN "0000000100100101" =>
						DD(2, 77) <= packet_in;
						counter <= "0000000100100110";
						WHEN "0000000100100110" =>
						DD(2, 78) <= packet_in;
						counter <= "0000000100100111";
						WHEN "0000000100100111" =>
						DD(2, 79) <= packet_in;
						counter <= "0000000100101000";
						WHEN "0000000100101000" =>
						DD(2, 80) <= packet_in;
						counter <= "0000000100101001";
						WHEN "0000000100101001" =>
						DD(2, 81) <= packet_in;
						counter <= "0000000100101010";
						WHEN "0000000100101010" =>
						DD(2, 82) <= packet_in;
						counter <= "0000000100101011";
						WHEN "0000000100101011" =>
						DD(2, 83) <= packet_in;
						counter <= "0000000100101100";
						WHEN "0000000100101100" =>
						DD(2, 84) <= packet_in;
						counter <= "0000000100101101";
						WHEN "0000000100101101" =>
						DD(2, 85) <= packet_in;
						counter <= "0000000100101110";
						WHEN "0000000100101110" =>
						DD(2, 86) <= packet_in;
						counter <= "0000000100101111";
						WHEN "0000000100101111" =>
						DD(2, 87) <= packet_in;
						counter <= "0000000100110000";
						WHEN "0000000100110000" =>
						DD(2, 88) <= packet_in;
						counter <= "0000000100110001";
						WHEN "0000000100110001" =>
						DD(2, 89) <= packet_in;
						counter <= "0000000100110010";
						WHEN "0000000100110010" =>
						DD(2, 90) <= packet_in;
						counter <= "0000000100110011";
						WHEN "0000000100110011" =>
						DD(2, 91) <= packet_in;
						counter <= "0000000100110100";
						WHEN "0000000100110100" =>
						DD(3, 0) <= packet_in;
						counter <= "0000000100110101";
						WHEN "0000000100110101" =>
						DD(3, 1) <= packet_in;
						counter <= "0000000100110110";
						WHEN "0000000100110110" =>
						DD(3, 2) <= packet_in;
						counter <= "0000000100110111";
						WHEN "0000000100110111" =>
						DD(3, 3) <= packet_in;
						counter <= "0000000100111000";
						WHEN "0000000100111000" =>
						DD(3, 4) <= packet_in;
						counter <= "0000000100111001";
						WHEN "0000000100111001" =>
						DD(3, 5) <= packet_in;
						counter <= "0000000100111010";
						WHEN "0000000100111010" =>
						DD(3, 6) <= packet_in;
						counter <= "0000000100111011";
						WHEN "0000000100111011" =>
						DD(3, 7) <= packet_in;
						counter <= "0000000100111100";
						WHEN "0000000100111100" =>
						DD(3, 8) <= packet_in;
						counter <= "0000000100111101";
						WHEN "0000000100111101" =>
						DD(3, 9) <= packet_in;
						counter <= "0000000100111110";
						WHEN "0000000100111110" =>
						DD(3, 10) <= packet_in;
						counter <= "0000000100111111";
						WHEN "0000000100111111" =>
						DD(3, 11) <= packet_in;
						counter <= "0000000101000000";
						WHEN "0000000101000000" =>
						DD(3, 12) <= packet_in;
						counter <= "0000000101000001";
						WHEN "0000000101000001" =>
						DD(3, 13) <= packet_in;
						counter <= "0000000101000010";
						WHEN "0000000101000010" =>
						DD(3, 14) <= packet_in;
						counter <= "0000000101000011";
						WHEN "0000000101000011" =>
						DD(3, 15) <= packet_in;
						counter <= "0000000101000100";
						WHEN "0000000101000100" =>
						DD(3, 16) <= packet_in;
						counter <= "0000000101000101";
						WHEN "0000000101000101" =>
						DD(3, 17) <= packet_in;
						counter <= "0000000101000110";
						WHEN "0000000101000110" =>
						DD(3, 18) <= packet_in;
						counter <= "0000000101000111";
						WHEN "0000000101000111" =>
						DD(3, 19) <= packet_in;
						counter <= "0000000101001000";
						WHEN "0000000101001000" =>
						DD(3, 20) <= packet_in;
						counter <= "0000000101001001";
						WHEN "0000000101001001" =>
						DD(3, 21) <= packet_in;
						counter <= "0000000101001010";
						WHEN "0000000101001010" =>
						DD(3, 22) <= packet_in;
						counter <= "0000000101001011";
						WHEN "0000000101001011" =>
						DD(3, 23) <= packet_in;
						counter <= "0000000101001100";
						WHEN "0000000101001100" =>
						DD(3, 24) <= packet_in;
						counter <= "0000000101001101";
						WHEN "0000000101001101" =>
						DD(3, 25) <= packet_in;
						counter <= "0000000101001110";
						WHEN "0000000101001110" =>
						DD(3, 26) <= packet_in;
						counter <= "0000000101001111";
						WHEN "0000000101001111" =>
						DD(3, 27) <= packet_in;
						counter <= "0000000101010000";
						WHEN "0000000101010000" =>
						DD(3, 28) <= packet_in;
						counter <= "0000000101010001";
						WHEN "0000000101010001" =>
						DD(3, 29) <= packet_in;
						counter <= "0000000101010010";
						WHEN "0000000101010010" =>
						DD(3, 30) <= packet_in;
						counter <= "0000000101010011";
						WHEN "0000000101010011" =>
						DD(3, 31) <= packet_in;
						counter <= "0000000101010100";
						WHEN "0000000101010100" =>
						DD(3, 32) <= packet_in;
						counter <= "0000000101010101";
						WHEN "0000000101010101" =>
						DD(3, 33) <= packet_in;
						counter <= "0000000101010110";
						WHEN "0000000101010110" =>
						DD(3, 34) <= packet_in;
						counter <= "0000000101010111";
						WHEN "0000000101010111" =>
						DD(3, 35) <= packet_in;
						counter <= "0000000101011000";
						WHEN "0000000101011000" =>
						DD(3, 36) <= packet_in;
						counter <= "0000000101011001";
						WHEN "0000000101011001" =>
						DD(3, 37) <= packet_in;
						counter <= "0000000101011010";
						WHEN "0000000101011010" =>
						DD(3, 38) <= packet_in;
						counter <= "0000000101011011";
						WHEN "0000000101011011" =>
						DD(3, 39) <= packet_in;
						counter <= "0000000101011100";
						WHEN "0000000101011100" =>
						DD(3, 40) <= packet_in;
						counter <= "0000000101011101";
						WHEN "0000000101011101" =>
						DD(3, 41) <= packet_in;
						counter <= "0000000101011110";
						WHEN "0000000101011110" =>
						DD(3, 42) <= packet_in;
						counter <= "0000000101011111";
						WHEN "0000000101011111" =>
						DD(3, 43) <= packet_in;
						counter <= "0000000101100000";
						WHEN "0000000101100000" =>
						DD(3, 44) <= packet_in;
						counter <= "0000000101100001";
						WHEN "0000000101100001" =>
						DD(3, 45) <= packet_in;
						counter <= "0000000101100010";
						WHEN "0000000101100010" =>
						DD(3, 46) <= packet_in;
						counter <= "0000000101100011";
						WHEN "0000000101100011" =>
						DD(3, 47) <= packet_in;
						counter <= "0000000101100100";
						WHEN "0000000101100100" =>
						DD(3, 48) <= packet_in;
						counter <= "0000000101100101";
						WHEN "0000000101100101" =>
						DD(3, 49) <= packet_in;
						counter <= "0000000101100110";
						WHEN "0000000101100110" =>
						DD(3, 50) <= packet_in;
						counter <= "0000000101100111";
						WHEN "0000000101100111" =>
						DD(3, 51) <= packet_in;
						counter <= "0000000101101000";
						WHEN "0000000101101000" =>
						DD(3, 52) <= packet_in;
						counter <= "0000000101101001";
						WHEN "0000000101101001" =>
						DD(3, 53) <= packet_in;
						counter <= "0000000101101010";
						WHEN "0000000101101010" =>
						DD(3, 54) <= packet_in;
						counter <= "0000000101101011";
						WHEN "0000000101101011" =>
						DD(3, 55) <= packet_in;
						counter <= "0000000101101100";
						WHEN "0000000101101100" =>
						DD(3, 56) <= packet_in;
						counter <= "0000000101101101";
						WHEN "0000000101101101" =>
						DD(3, 57) <= packet_in;
						counter <= "0000000101101110";
						WHEN "0000000101101110" =>
						DD(3, 58) <= packet_in;
						counter <= "0000000101101111";
						WHEN "0000000101101111" =>
						DD(3, 59) <= packet_in;
						counter <= "0000000101110000";
						WHEN "0000000101110000" =>
						DD(3, 60) <= packet_in;
						counter <= "0000000101110001";
						WHEN "0000000101110001" =>
						DD(3, 61) <= packet_in;
						counter <= "0000000101110010";
						WHEN "0000000101110010" =>
						DD(3, 62) <= packet_in;
						counter <= "0000000101110011";
						WHEN "0000000101110011" =>
						DD(3, 63) <= packet_in;
						counter <= "0000000101110100";
						WHEN "0000000101110100" =>
						DD(3, 64) <= packet_in;
						counter <= "0000000101110101";
						WHEN "0000000101110101" =>
						DD(3, 65) <= packet_in;
						counter <= "0000000101110110";
						WHEN "0000000101110110" =>
						DD(3, 66) <= packet_in;
						counter <= "0000000101110111";
						WHEN "0000000101110111" =>
						DD(3, 67) <= packet_in;
						counter <= "0000000101111000";
						WHEN "0000000101111000" =>
						DD(3, 68) <= packet_in;
						counter <= "0000000101111001";
						WHEN "0000000101111001" =>
						DD(3, 69) <= packet_in;
						counter <= "0000000101111010";
						WHEN "0000000101111010" =>
						DD(3, 70) <= packet_in;
						counter <= "0000000101111011";
						WHEN "0000000101111011" =>
						DD(3, 71) <= packet_in;
						counter <= "0000000101111100";
						WHEN "0000000101111100" =>
						DD(3, 72) <= packet_in;
						counter <= "0000000101111101";
						WHEN "0000000101111101" =>
						DD(3, 73) <= packet_in;
						counter <= "0000000101111110";
						WHEN "0000000101111110" =>
						DD(3, 74) <= packet_in;
						counter <= "0000000101111111";
						WHEN "0000000101111111" =>
						DD(3, 75) <= packet_in;
						counter <= "0000000110000000";
						WHEN "0000000110000000" =>
						DD(3, 76) <= packet_in;
						counter <= "0000000110000001";
						WHEN "0000000110000001" =>
						DD(3, 77) <= packet_in;
						counter <= "0000000110000010";
						WHEN "0000000110000010" =>
						DD(3, 78) <= packet_in;
						counter <= "0000000110000011";
						WHEN "0000000110000011" =>
						DD(3, 79) <= packet_in;
						counter <= "0000000110000100";
						WHEN "0000000110000100" =>
						DD(3, 80) <= packet_in;
						counter <= "0000000110000101";
						WHEN "0000000110000101" =>
						DD(3, 81) <= packet_in;
						counter <= "0000000110000110";
						WHEN "0000000110000110" =>
						DD(3, 82) <= packet_in;
						counter <= "0000000110000111";
						WHEN "0000000110000111" =>
						DD(3, 83) <= packet_in;
						counter <= "0000000110001000";
						WHEN "0000000110001000" =>
						DD(3, 84) <= packet_in;
						counter <= "0000000110001001";
						WHEN "0000000110001001" =>
						DD(3, 85) <= packet_in;
						counter <= "0000000110001010";
						WHEN "0000000110001010" =>
						DD(3, 86) <= packet_in;
						counter <= "0000000110001011";
						WHEN "0000000110001011" =>
						DD(3, 87) <= packet_in;
						counter <= "0000000110001100";
						WHEN "0000000110001100" =>
						DD(3, 88) <= packet_in;
						counter <= "0000000110001101";
						WHEN "0000000110001101" =>
						DD(3, 89) <= packet_in;
						counter <= "0000000110001110";
						WHEN "0000000110001110" =>
						DD(3, 90) <= packet_in;
						counter <= "0000000110001111";
						WHEN "0000000110001111" =>
						DD(3, 91) <= packet_in;
						counter <= "0000000110010000";
						WHEN "0000000110010000" =>
						DD(4, 0) <= packet_in;
						counter <= "0000000110010001";
						WHEN "0000000110010001" =>
						DD(4, 1) <= packet_in;
						counter <= "0000000110010010";
						WHEN "0000000110010010" =>
						DD(4, 2) <= packet_in;
						counter <= "0000000110010011";
						WHEN "0000000110010011" =>
						DD(4, 3) <= packet_in;
						counter <= "0000000110010100";
						WHEN "0000000110010100" =>
						DD(4, 4) <= packet_in;
						counter <= "0000000110010101";
						WHEN "0000000110010101" =>
						DD(4, 5) <= packet_in;
						counter <= "0000000110010110";
						WHEN "0000000110010110" =>
						DD(4, 6) <= packet_in;
						counter <= "0000000110010111";
						WHEN "0000000110010111" =>
						DD(4, 7) <= packet_in;
						counter <= "0000000110011000";
						WHEN "0000000110011000" =>
						DD(4, 8) <= packet_in;
						counter <= "0000000110011001";
						WHEN "0000000110011001" =>
						DD(4, 9) <= packet_in;
						counter <= "0000000110011010";
						WHEN "0000000110011010" =>
						DD(4, 10) <= packet_in;
						counter <= "0000000110011011";
						WHEN "0000000110011011" =>
						DD(4, 11) <= packet_in;
						counter <= "0000000110011100";
						WHEN "0000000110011100" =>
						DD(4, 12) <= packet_in;
						counter <= "0000000110011101";
						WHEN "0000000110011101" =>
						DD(4, 13) <= packet_in;
						counter <= "0000000110011110";
						WHEN "0000000110011110" =>
						DD(4, 14) <= packet_in;
						counter <= "0000000110011111";
						WHEN "0000000110011111" =>
						DD(4, 15) <= packet_in;
						counter <= "0000000110100000";
						WHEN "0000000110100000" =>
						DD(4, 16) <= packet_in;
						counter <= "0000000110100001";
						WHEN "0000000110100001" =>
						DD(4, 17) <= packet_in;
						counter <= "0000000110100010";
						WHEN "0000000110100010" =>
						DD(4, 18) <= packet_in;
						counter <= "0000000110100011";
						WHEN "0000000110100011" =>
						DD(4, 19) <= packet_in;
						counter <= "0000000110100100";
						WHEN "0000000110100100" =>
						DD(4, 20) <= packet_in;
						counter <= "0000000110100101";
						WHEN "0000000110100101" =>
						DD(4, 21) <= packet_in;
						counter <= "0000000110100110";
						WHEN "0000000110100110" =>
						DD(4, 22) <= packet_in;
						counter <= "0000000110100111";
						WHEN "0000000110100111" =>
						DD(4, 23) <= packet_in;
						counter <= "0000000110101000";
						WHEN "0000000110101000" =>
						DD(4, 24) <= packet_in;
						counter <= "0000000110101001";
						WHEN "0000000110101001" =>
						DD(4, 25) <= packet_in;
						counter <= "0000000110101010";
						WHEN "0000000110101010" =>
						DD(4, 26) <= packet_in;
						counter <= "0000000110101011";
						WHEN "0000000110101011" =>
						DD(4, 27) <= packet_in;
						counter <= "0000000110101100";
						WHEN "0000000110101100" =>
						DD(4, 28) <= packet_in;
						counter <= "0000000110101101";
						WHEN "0000000110101101" =>
						DD(4, 29) <= packet_in;
						counter <= "0000000110101110";
						WHEN "0000000110101110" =>
						DD(4, 30) <= packet_in;
						counter <= "0000000110101111";
						WHEN "0000000110101111" =>
						DD(4, 31) <= packet_in;
						counter <= "0000000110110000";
						WHEN "0000000110110000" =>
						DD(4, 32) <= packet_in;
						counter <= "0000000110110001";
						WHEN "0000000110110001" =>
						DD(4, 33) <= packet_in;
						counter <= "0000000110110010";
						WHEN "0000000110110010" =>
						DD(4, 34) <= packet_in;
						counter <= "0000000110110011";
						WHEN "0000000110110011" =>
						DD(4, 35) <= packet_in;
						counter <= "0000000110110100";
						WHEN "0000000110110100" =>
						DD(4, 36) <= packet_in;
						counter <= "0000000110110101";
						WHEN "0000000110110101" =>
						DD(4, 37) <= packet_in;
						counter <= "0000000110110110";
						WHEN "0000000110110110" =>
						DD(4, 38) <= packet_in;
						counter <= "0000000110110111";
						WHEN "0000000110110111" =>
						DD(4, 39) <= packet_in;
						counter <= "0000000110111000";
						WHEN "0000000110111000" =>
						DD(4, 40) <= packet_in;
						counter <= "0000000110111001";
						WHEN "0000000110111001" =>
						DD(4, 41) <= packet_in;
						counter <= "0000000110111010";
						WHEN "0000000110111010" =>
						DD(4, 42) <= packet_in;
						counter <= "0000000110111011";
						WHEN "0000000110111011" =>
						DD(4, 43) <= packet_in;
						counter <= "0000000110111100";
						WHEN "0000000110111100" =>
						DD(4, 44) <= packet_in;
						counter <= "0000000110111101";
						WHEN "0000000110111101" =>
						DD(4, 45) <= packet_in;
						counter <= "0000000110111110";
						WHEN "0000000110111110" =>
						DD(4, 46) <= packet_in;
						counter <= "0000000110111111";
						WHEN "0000000110111111" =>
						DD(4, 47) <= packet_in;
						counter <= "0000000111000000";
						WHEN "0000000111000000" =>
						DD(4, 48) <= packet_in;
						counter <= "0000000111000001";
						WHEN "0000000111000001" =>
						DD(4, 49) <= packet_in;
						counter <= "0000000111000010";
						WHEN "0000000111000010" =>
						DD(4, 50) <= packet_in;
						counter <= "0000000111000011";
						WHEN "0000000111000011" =>
						DD(4, 51) <= packet_in;
						counter <= "0000000111000100";
						WHEN "0000000111000100" =>
						DD(4, 52) <= packet_in;
						counter <= "0000000111000101";
						WHEN "0000000111000101" =>
						DD(4, 53) <= packet_in;
						counter <= "0000000111000110";
						WHEN "0000000111000110" =>
						DD(4, 54) <= packet_in;
						counter <= "0000000111000111";
						WHEN "0000000111000111" =>
						DD(4, 55) <= packet_in;
						counter <= "0000000111001000";
						WHEN "0000000111001000" =>
						DD(4, 56) <= packet_in;
						counter <= "0000000111001001";
						WHEN "0000000111001001" =>
						DD(4, 57) <= packet_in;
						counter <= "0000000111001010";
						WHEN "0000000111001010" =>
						DD(4, 58) <= packet_in;
						counter <= "0000000111001011";
						WHEN "0000000111001011" =>
						DD(4, 59) <= packet_in;
						counter <= "0000000111001100";
						WHEN "0000000111001100" =>
						DD(4, 60) <= packet_in;
						counter <= "0000000111001101";
						WHEN "0000000111001101" =>
						DD(4, 61) <= packet_in;
						counter <= "0000000111001110";
						WHEN "0000000111001110" =>
						DD(4, 62) <= packet_in;
						counter <= "0000000111001111";
						WHEN "0000000111001111" =>
						DD(4, 63) <= packet_in;
						counter <= "0000000111010000";
						WHEN "0000000111010000" =>
						DD(4, 64) <= packet_in;
						counter <= "0000000111010001";
						WHEN "0000000111010001" =>
						DD(4, 65) <= packet_in;
						counter <= "0000000111010010";
						WHEN "0000000111010010" =>
						DD(4, 66) <= packet_in;
						counter <= "0000000111010011";
						WHEN "0000000111010011" =>
						DD(4, 67) <= packet_in;
						counter <= "0000000111010100";
						WHEN "0000000111010100" =>
						DD(4, 68) <= packet_in;
						counter <= "0000000111010101";
						WHEN "0000000111010101" =>
						DD(4, 69) <= packet_in;
						counter <= "0000000111010110";
						WHEN "0000000111010110" =>
						DD(4, 70) <= packet_in;
						counter <= "0000000111010111";
						WHEN "0000000111010111" =>
						DD(4, 71) <= packet_in;
						counter <= "0000000111011000";
						WHEN "0000000111011000" =>
						DD(4, 72) <= packet_in;
						counter <= "0000000111011001";
						WHEN "0000000111011001" =>
						DD(4, 73) <= packet_in;
						counter <= "0000000111011010";
						WHEN "0000000111011010" =>
						DD(4, 74) <= packet_in;
						counter <= "0000000111011011";
						WHEN "0000000111011011" =>
						DD(4, 75) <= packet_in;
						counter <= "0000000111011100";
						WHEN "0000000111011100" =>
						DD(4, 76) <= packet_in;
						counter <= "0000000111011101";
						WHEN "0000000111011101" =>
						DD(4, 77) <= packet_in;
						counter <= "0000000111011110";
						WHEN "0000000111011110" =>
						DD(4, 78) <= packet_in;
						counter <= "0000000111011111";
						WHEN "0000000111011111" =>
						DD(4, 79) <= packet_in;
						counter <= "0000000111100000";
						WHEN "0000000111100000" =>
						DD(4, 80) <= packet_in;
						counter <= "0000000111100001";
						WHEN "0000000111100001" =>
						DD(4, 81) <= packet_in;
						counter <= "0000000111100010";
						WHEN "0000000111100010" =>
						DD(4, 82) <= packet_in;
						counter <= "0000000111100011";
						WHEN "0000000111100011" =>
						DD(4, 83) <= packet_in;
						counter <= "0000000111100100";
						WHEN "0000000111100100" =>
						DD(4, 84) <= packet_in;
						counter <= "0000000111100101";
						WHEN "0000000111100101" =>
						DD(4, 85) <= packet_in;
						counter <= "0000000111100110";
						WHEN "0000000111100110" =>
						DD(4, 86) <= packet_in;
						counter <= "0000000111100111";
						WHEN "0000000111100111" =>
						DD(4, 87) <= packet_in;
						counter <= "0000000111101000";
						WHEN "0000000111101000" =>
						DD(4, 88) <= packet_in;
						counter <= "0000000111101001";
						WHEN "0000000111101001" =>
						DD(4, 89) <= packet_in;
						counter <= "0000000111101010";
						WHEN "0000000111101010" =>
						DD(4, 90) <= packet_in;
						counter <= "0000000111101011";
						WHEN "0000000111101011" =>
						DD(4, 91) <= packet_in;
						counter <= "0000000111101100";
						WHEN "0000000111101100" =>
						DD(5, 0) <= packet_in;
						counter <= "0000000111101101";
						WHEN "0000000111101101" =>
						DD(5, 1) <= packet_in;
						counter <= "0000000111101110";
						WHEN "0000000111101110" =>
						DD(5, 2) <= packet_in;
						counter <= "0000000111101111";
						WHEN "0000000111101111" =>
						DD(5, 3) <= packet_in;
						counter <= "0000000111110000";
						WHEN "0000000111110000" =>
						DD(5, 4) <= packet_in;
						counter <= "0000000111110001";
						WHEN "0000000111110001" =>
						DD(5, 5) <= packet_in;
						counter <= "0000000111110010";
						WHEN "0000000111110010" =>
						DD(5, 6) <= packet_in;
						counter <= "0000000111110011";
						WHEN "0000000111110011" =>
						DD(5, 7) <= packet_in;
						counter <= "0000000111110100";
						WHEN "0000000111110100" =>
						DD(5, 8) <= packet_in;
						counter <= "0000000111110101";
						WHEN "0000000111110101" =>
						DD(5, 9) <= packet_in;
						counter <= "0000000111110110";
						WHEN "0000000111110110" =>
						DD(5, 10) <= packet_in;
						counter <= "0000000111110111";
						WHEN "0000000111110111" =>
						DD(5, 11) <= packet_in;
						counter <= "0000000111111000";
						WHEN "0000000111111000" =>
						DD(5, 12) <= packet_in;
						counter <= "0000000111111001";
						WHEN "0000000111111001" =>
						DD(5, 13) <= packet_in;
						counter <= "0000000111111010";
						WHEN "0000000111111010" =>
						DD(5, 14) <= packet_in;
						counter <= "0000000111111011";
						WHEN "0000000111111011" =>
						DD(5, 15) <= packet_in;
						counter <= "0000000111111100";
						WHEN "0000000111111100" =>
						DD(5, 16) <= packet_in;
						counter <= "0000000111111101";
						WHEN "0000000111111101" =>
						DD(5, 17) <= packet_in;
						counter <= "0000000111111110";
						WHEN "0000000111111110" =>
						DD(5, 18) <= packet_in;
						counter <= "0000000111111111";
						WHEN "0000000111111111" =>
						DD(5, 19) <= packet_in;
						counter <= "0000001000000000";
						WHEN "0000001000000000" =>
						DD(5, 20) <= packet_in;
						counter <= "0000001000000001";
						WHEN "0000001000000001" =>
						DD(5, 21) <= packet_in;
						counter <= "0000001000000010";
						WHEN "0000001000000010" =>
						DD(5, 22) <= packet_in;
						counter <= "0000001000000011";
						WHEN "0000001000000011" =>
						DD(5, 23) <= packet_in;
						counter <= "0000001000000100";
						WHEN "0000001000000100" =>
						DD(5, 24) <= packet_in;
						counter <= "0000001000000101";
						WHEN "0000001000000101" =>
						DD(5, 25) <= packet_in;
						counter <= "0000001000000110";
						WHEN "0000001000000110" =>
						DD(5, 26) <= packet_in;
						counter <= "0000001000000111";
						WHEN "0000001000000111" =>
						DD(5, 27) <= packet_in;
						counter <= "0000001000001000";
						WHEN "0000001000001000" =>
						DD(5, 28) <= packet_in;
						counter <= "0000001000001001";
						WHEN "0000001000001001" =>
						DD(5, 29) <= packet_in;
						counter <= "0000001000001010";
						WHEN "0000001000001010" =>
						DD(5, 30) <= packet_in;
						counter <= "0000001000001011";
						WHEN "0000001000001011" =>
						DD(5, 31) <= packet_in;
						counter <= "0000001000001100";
						WHEN "0000001000001100" =>
						DD(5, 32) <= packet_in;
						counter <= "0000001000001101";
						WHEN "0000001000001101" =>
						DD(5, 33) <= packet_in;
						counter <= "0000001000001110";
						WHEN "0000001000001110" =>
						DD(5, 34) <= packet_in;
						counter <= "0000001000001111";
						WHEN "0000001000001111" =>
						DD(5, 35) <= packet_in;
						counter <= "0000001000010000";
						WHEN "0000001000010000" =>
						DD(5, 36) <= packet_in;
						counter <= "0000001000010001";
						WHEN "0000001000010001" =>
						DD(5, 37) <= packet_in;
						counter <= "0000001000010010";
						WHEN "0000001000010010" =>
						DD(5, 38) <= packet_in;
						counter <= "0000001000010011";
						WHEN "0000001000010011" =>
						DD(5, 39) <= packet_in;
						counter <= "0000001000010100";
						WHEN "0000001000010100" =>
						DD(5, 40) <= packet_in;
						counter <= "0000001000010101";
						WHEN "0000001000010101" =>
						DD(5, 41) <= packet_in;
						counter <= "0000001000010110";
						WHEN "0000001000010110" =>
						DD(5, 42) <= packet_in;
						counter <= "0000001000010111";
						WHEN "0000001000010111" =>
						DD(5, 43) <= packet_in;
						counter <= "0000001000011000";
						WHEN "0000001000011000" =>
						DD(5, 44) <= packet_in;
						counter <= "0000001000011001";
						WHEN "0000001000011001" =>
						DD(5, 45) <= packet_in;
						counter <= "0000001000011010";
						WHEN "0000001000011010" =>
						DD(5, 46) <= packet_in;
						counter <= "0000001000011011";
						WHEN "0000001000011011" =>
						DD(5, 47) <= packet_in;
						counter <= "0000001000011100";
						WHEN "0000001000011100" =>
						DD(5, 48) <= packet_in;
						counter <= "0000001000011101";
						WHEN "0000001000011101" =>
						DD(5, 49) <= packet_in;
						counter <= "0000001000011110";
						WHEN "0000001000011110" =>
						DD(5, 50) <= packet_in;
						counter <= "0000001000011111";
						WHEN "0000001000011111" =>
						DD(5, 51) <= packet_in;
						counter <= "0000001000100000";
						WHEN "0000001000100000" =>
						DD(5, 52) <= packet_in;
						counter <= "0000001000100001";
						WHEN "0000001000100001" =>
						DD(5, 53) <= packet_in;
						counter <= "0000001000100010";
						WHEN "0000001000100010" =>
						DD(5, 54) <= packet_in;
						counter <= "0000001000100011";
						WHEN "0000001000100011" =>
						DD(5, 55) <= packet_in;
						counter <= "0000001000100100";
						WHEN "0000001000100100" =>
						DD(5, 56) <= packet_in;
						counter <= "0000001000100101";
						WHEN "0000001000100101" =>
						DD(5, 57) <= packet_in;
						counter <= "0000001000100110";
						WHEN "0000001000100110" =>
						DD(5, 58) <= packet_in;
						counter <= "0000001000100111";
						WHEN "0000001000100111" =>
						DD(5, 59) <= packet_in;
						counter <= "0000001000101000";
						WHEN "0000001000101000" =>
						DD(5, 60) <= packet_in;
						counter <= "0000001000101001";
						WHEN "0000001000101001" =>
						DD(5, 61) <= packet_in;
						counter <= "0000001000101010";
						WHEN "0000001000101010" =>
						DD(5, 62) <= packet_in;
						counter <= "0000001000101011";
						WHEN "0000001000101011" =>
						DD(5, 63) <= packet_in;
						counter <= "0000001000101100";
						WHEN "0000001000101100" =>
						DD(5, 64) <= packet_in;
						counter <= "0000001000101101";
						WHEN "0000001000101101" =>
						DD(5, 65) <= packet_in;
						counter <= "0000001000101110";
						WHEN "0000001000101110" =>
						DD(5, 66) <= packet_in;
						counter <= "0000001000101111";
						WHEN "0000001000101111" =>
						DD(5, 67) <= packet_in;
						counter <= "0000001000110000";
						WHEN "0000001000110000" =>
						DD(5, 68) <= packet_in;
						counter <= "0000001000110001";
						WHEN "0000001000110001" =>
						DD(5, 69) <= packet_in;
						counter <= "0000001000110010";
						WHEN "0000001000110010" =>
						DD(5, 70) <= packet_in;
						counter <= "0000001000110011";
						WHEN "0000001000110011" =>
						DD(5, 71) <= packet_in;
						counter <= "0000001000110100";
						WHEN "0000001000110100" =>
						DD(5, 72) <= packet_in;
						counter <= "0000001000110101";
						WHEN "0000001000110101" =>
						DD(5, 73) <= packet_in;
						counter <= "0000001000110110";
						WHEN "0000001000110110" =>
						DD(5, 74) <= packet_in;
						counter <= "0000001000110111";
						WHEN "0000001000110111" =>
						DD(5, 75) <= packet_in;
						counter <= "0000001000111000";
						WHEN "0000001000111000" =>
						DD(5, 76) <= packet_in;
						counter <= "0000001000111001";
						WHEN "0000001000111001" =>
						DD(5, 77) <= packet_in;
						counter <= "0000001000111010";
						WHEN "0000001000111010" =>
						DD(5, 78) <= packet_in;
						counter <= "0000001000111011";
						WHEN "0000001000111011" =>
						DD(5, 79) <= packet_in;
						counter <= "0000001000111100";
						WHEN "0000001000111100" =>
						DD(5, 80) <= packet_in;
						counter <= "0000001000111101";
						WHEN "0000001000111101" =>
						DD(5, 81) <= packet_in;
						counter <= "0000001000111110";
						WHEN "0000001000111110" =>
						DD(5, 82) <= packet_in;
						counter <= "0000001000111111";
						WHEN "0000001000111111" =>
						DD(5, 83) <= packet_in;
						counter <= "0000001001000000";
						WHEN "0000001001000000" =>
						DD(5, 84) <= packet_in;
						counter <= "0000001001000001";
						WHEN "0000001001000001" =>
						DD(5, 85) <= packet_in;
						counter <= "0000001001000010";
						WHEN "0000001001000010" =>
						DD(5, 86) <= packet_in;
						counter <= "0000001001000011";
						WHEN "0000001001000011" =>
						DD(5, 87) <= packet_in;
						counter <= "0000001001000100";
						WHEN "0000001001000100" =>
						DD(5, 88) <= packet_in;
						counter <= "0000001001000101";
						WHEN "0000001001000101" =>
						DD(5, 89) <= packet_in;
						counter <= "0000001001000110";
						WHEN "0000001001000110" =>
						DD(5, 90) <= packet_in;
						counter <= "0000001001000111";
						WHEN "0000001001000111" =>
						DD(5, 91) <= packet_in;
						counter <= "0000001001001000";
						WHEN "0000001001001000" =>
						DD(6, 0) <= packet_in;
						counter <= "0000001001001001";
						WHEN "0000001001001001" =>
						DD(6, 1) <= packet_in;
						counter <= "0000001001001010";
						WHEN "0000001001001010" =>
						DD(6, 2) <= packet_in;
						counter <= "0000001001001011";
						WHEN "0000001001001011" =>
						DD(6, 3) <= packet_in;
						counter <= "0000001001001100";
						WHEN "0000001001001100" =>
						DD(6, 4) <= packet_in;
						counter <= "0000001001001101";
						WHEN "0000001001001101" =>
						DD(6, 5) <= packet_in;
						counter <= "0000001001001110";
						WHEN "0000001001001110" =>
						DD(6, 6) <= packet_in;
						counter <= "0000001001001111";
						WHEN "0000001001001111" =>
						DD(6, 7) <= packet_in;
						counter <= "0000001001010000";
						WHEN "0000001001010000" =>
						DD(6, 8) <= packet_in;
						counter <= "0000001001010001";
						WHEN "0000001001010001" =>
						DD(6, 9) <= packet_in;
						counter <= "0000001001010010";
						WHEN "0000001001010010" =>
						DD(6, 10) <= packet_in;
						counter <= "0000001001010011";
						WHEN "0000001001010011" =>
						DD(6, 11) <= packet_in;
						counter <= "0000001001010100";
						WHEN "0000001001010100" =>
						DD(6, 12) <= packet_in;
						counter <= "0000001001010101";
						WHEN "0000001001010101" =>
						DD(6, 13) <= packet_in;
						counter <= "0000001001010110";
						WHEN "0000001001010110" =>
						DD(6, 14) <= packet_in;
						counter <= "0000001001010111";
						WHEN "0000001001010111" =>
						DD(6, 15) <= packet_in;
						counter <= "0000001001011000";
						WHEN "0000001001011000" =>
						DD(6, 16) <= packet_in;
						counter <= "0000001001011001";
						WHEN "0000001001011001" =>
						DD(6, 17) <= packet_in;
						counter <= "0000001001011010";
						WHEN "0000001001011010" =>
						DD(6, 18) <= packet_in;
						counter <= "0000001001011011";
						WHEN "0000001001011011" =>
						DD(6, 19) <= packet_in;
						counter <= "0000001001011100";
						WHEN "0000001001011100" =>
						DD(6, 20) <= packet_in;
						counter <= "0000001001011101";
						WHEN "0000001001011101" =>
						DD(6, 21) <= packet_in;
						counter <= "0000001001011110";
						WHEN "0000001001011110" =>
						DD(6, 22) <= packet_in;
						counter <= "0000001001011111";
						WHEN "0000001001011111" =>
						DD(6, 23) <= packet_in;
						counter <= "0000001001100000";
						WHEN "0000001001100000" =>
						DD(6, 24) <= packet_in;
						counter <= "0000001001100001";
						WHEN "0000001001100001" =>
						DD(6, 25) <= packet_in;
						counter <= "0000001001100010";
						WHEN "0000001001100010" =>
						DD(6, 26) <= packet_in;
						counter <= "0000001001100011";
						WHEN "0000001001100011" =>
						DD(6, 27) <= packet_in;
						counter <= "0000001001100100";
						WHEN "0000001001100100" =>
						DD(6, 28) <= packet_in;
						counter <= "0000001001100101";
						WHEN "0000001001100101" =>
						DD(6, 29) <= packet_in;
						counter <= "0000001001100110";
						WHEN "0000001001100110" =>
						DD(6, 30) <= packet_in;
						counter <= "0000001001100111";
						WHEN "0000001001100111" =>
						DD(6, 31) <= packet_in;
						counter <= "0000001001101000";
						WHEN "0000001001101000" =>
						DD(6, 32) <= packet_in;
						counter <= "0000001001101001";
						WHEN "0000001001101001" =>
						DD(6, 33) <= packet_in;
						counter <= "0000001001101010";
						WHEN "0000001001101010" =>
						DD(6, 34) <= packet_in;
						counter <= "0000001001101011";
						WHEN "0000001001101011" =>
						DD(6, 35) <= packet_in;
						counter <= "0000001001101100";
						WHEN "0000001001101100" =>
						DD(6, 36) <= packet_in;
						counter <= "0000001001101101";
						WHEN "0000001001101101" =>
						DD(6, 37) <= packet_in;
						counter <= "0000001001101110";
						WHEN "0000001001101110" =>
						DD(6, 38) <= packet_in;
						counter <= "0000001001101111";
						WHEN "0000001001101111" =>
						DD(6, 39) <= packet_in;
						counter <= "0000001001110000";
						WHEN "0000001001110000" =>
						DD(6, 40) <= packet_in;
						counter <= "0000001001110001";
						WHEN "0000001001110001" =>
						DD(6, 41) <= packet_in;
						counter <= "0000001001110010";
						WHEN "0000001001110010" =>
						DD(6, 42) <= packet_in;
						counter <= "0000001001110011";
						WHEN "0000001001110011" =>
						DD(6, 43) <= packet_in;
						counter <= "0000001001110100";
						WHEN "0000001001110100" =>
						DD(6, 44) <= packet_in;
						counter <= "0000001001110101";
						WHEN "0000001001110101" =>
						DD(6, 45) <= packet_in;
						counter <= "0000001001110110";
						WHEN "0000001001110110" =>
						DD(6, 46) <= packet_in;
						counter <= "0000001001110111";
						WHEN "0000001001110111" =>
						DD(6, 47) <= packet_in;
						counter <= "0000001001111000";
						WHEN "0000001001111000" =>
						DD(6, 48) <= packet_in;
						counter <= "0000001001111001";
						WHEN "0000001001111001" =>
						DD(6, 49) <= packet_in;
						counter <= "0000001001111010";
						WHEN "0000001001111010" =>
						DD(6, 50) <= packet_in;
						counter <= "0000001001111011";
						WHEN "0000001001111011" =>
						DD(6, 51) <= packet_in;
						counter <= "0000001001111100";
						WHEN "0000001001111100" =>
						DD(6, 52) <= packet_in;
						counter <= "0000001001111101";
						WHEN "0000001001111101" =>
						DD(6, 53) <= packet_in;
						counter <= "0000001001111110";
						WHEN "0000001001111110" =>
						DD(6, 54) <= packet_in;
						counter <= "0000001001111111";
						WHEN "0000001001111111" =>
						DD(6, 55) <= packet_in;
						counter <= "0000001010000000";
						WHEN "0000001010000000" =>
						DD(6, 56) <= packet_in;
						counter <= "0000001010000001";
						WHEN "0000001010000001" =>
						DD(6, 57) <= packet_in;
						counter <= "0000001010000010";
						WHEN "0000001010000010" =>
						DD(6, 58) <= packet_in;
						counter <= "0000001010000011";
						WHEN "0000001010000011" =>
						DD(6, 59) <= packet_in;
						counter <= "0000001010000100";
						WHEN "0000001010000100" =>
						DD(6, 60) <= packet_in;
						counter <= "0000001010000101";
						WHEN "0000001010000101" =>
						DD(6, 61) <= packet_in;
						counter <= "0000001010000110";
						WHEN "0000001010000110" =>
						DD(6, 62) <= packet_in;
						counter <= "0000001010000111";
						WHEN "0000001010000111" =>
						DD(6, 63) <= packet_in;
						counter <= "0000001010001000";
						WHEN "0000001010001000" =>
						DD(6, 64) <= packet_in;
						counter <= "0000001010001001";
						WHEN "0000001010001001" =>
						DD(6, 65) <= packet_in;
						counter <= "0000001010001010";
						WHEN "0000001010001010" =>
						DD(6, 66) <= packet_in;
						counter <= "0000001010001011";
						WHEN "0000001010001011" =>
						DD(6, 67) <= packet_in;
						counter <= "0000001010001100";
						WHEN "0000001010001100" =>
						DD(6, 68) <= packet_in;
						counter <= "0000001010001101";
						WHEN "0000001010001101" =>
						DD(6, 69) <= packet_in;
						counter <= "0000001010001110";
						WHEN "0000001010001110" =>
						DD(6, 70) <= packet_in;
						counter <= "0000001010001111";
						WHEN "0000001010001111" =>
						DD(6, 71) <= packet_in;
						counter <= "0000001010010000";
						WHEN "0000001010010000" =>
						DD(6, 72) <= packet_in;
						counter <= "0000001010010001";
						WHEN "0000001010010001" =>
						DD(6, 73) <= packet_in;
						counter <= "0000001010010010";
						WHEN "0000001010010010" =>
						DD(6, 74) <= packet_in;
						counter <= "0000001010010011";
						WHEN "0000001010010011" =>
						DD(6, 75) <= packet_in;
						counter <= "0000001010010100";
						WHEN "0000001010010100" =>
						DD(6, 76) <= packet_in;
						counter <= "0000001010010101";
						WHEN "0000001010010101" =>
						DD(6, 77) <= packet_in;
						counter <= "0000001010010110";
						WHEN "0000001010010110" =>
						DD(6, 78) <= packet_in;
						counter <= "0000001010010111";
						WHEN "0000001010010111" =>
						DD(6, 79) <= packet_in;
						counter <= "0000001010011000";
						WHEN "0000001010011000" =>
						DD(6, 80) <= packet_in;
						counter <= "0000001010011001";
						WHEN "0000001010011001" =>
						DD(6, 81) <= packet_in;
						counter <= "0000001010011010";
						WHEN "0000001010011010" =>
						DD(6, 82) <= packet_in;
						counter <= "0000001010011011";
						WHEN "0000001010011011" =>
						DD(6, 83) <= packet_in;
						counter <= "0000001010011100";
						WHEN "0000001010011100" =>
						DD(6, 84) <= packet_in;
						counter <= "0000001010011101";
						WHEN "0000001010011101" =>
						DD(6, 85) <= packet_in;
						counter <= "0000001010011110";
						WHEN "0000001010011110" =>
						DD(6, 86) <= packet_in;
						counter <= "0000001010011111";
						WHEN "0000001010011111" =>
						DD(6, 87) <= packet_in;
						counter <= "0000001010100000";
						WHEN "0000001010100000" =>
						DD(6, 88) <= packet_in;
						counter <= "0000001010100001";
						WHEN "0000001010100001" =>
						DD(6, 89) <= packet_in;
						counter <= "0000001010100010";
						WHEN "0000001010100010" =>
						DD(6, 90) <= packet_in;
						counter <= "0000001010100011";
						WHEN "0000001010100011" =>
						DD(6, 91) <= packet_in;
						counter <= "0000001010100100";
						WHEN "0000001010100100" =>
						DD(7, 0) <= packet_in;
						counter <= "0000001010100101";
						WHEN "0000001010100101" =>
						DD(7, 1) <= packet_in;
						counter <= "0000001010100110";
						WHEN "0000001010100110" =>
						DD(7, 2) <= packet_in;
						counter <= "0000001010100111";
						WHEN "0000001010100111" =>
						DD(7, 3) <= packet_in;
						counter <= "0000001010101000";
						WHEN "0000001010101000" =>
						DD(7, 4) <= packet_in;
						counter <= "0000001010101001";
						WHEN "0000001010101001" =>
						DD(7, 5) <= packet_in;
						counter <= "0000001010101010";
						WHEN "0000001010101010" =>
						DD(7, 6) <= packet_in;
						counter <= "0000001010101011";
						WHEN "0000001010101011" =>
						DD(7, 7) <= packet_in;
						counter <= "0000001010101100";
						WHEN "0000001010101100" =>
						DD(7, 8) <= packet_in;
						counter <= "0000001010101101";
						WHEN "0000001010101101" =>
						DD(7, 9) <= packet_in;
						counter <= "0000001010101110";
						WHEN "0000001010101110" =>
						DD(7, 10) <= packet_in;
						counter <= "0000001010101111";
						WHEN "0000001010101111" =>
						DD(7, 11) <= packet_in;
						counter <= "0000001010110000";
						WHEN "0000001010110000" =>
						DD(7, 12) <= packet_in;
						counter <= "0000001010110001";
						WHEN "0000001010110001" =>
						DD(7, 13) <= packet_in;
						counter <= "0000001010110010";
						WHEN "0000001010110010" =>
						DD(7, 14) <= packet_in;
						counter <= "0000001010110011";
						WHEN "0000001010110011" =>
						DD(7, 15) <= packet_in;
						counter <= "0000001010110100";
						WHEN "0000001010110100" =>
						DD(7, 16) <= packet_in;
						counter <= "0000001010110101";
						WHEN "0000001010110101" =>
						DD(7, 17) <= packet_in;
						counter <= "0000001010110110";
						WHEN "0000001010110110" =>
						DD(7, 18) <= packet_in;
						counter <= "0000001010110111";
						WHEN "0000001010110111" =>
						DD(7, 19) <= packet_in;
						counter <= "0000001010111000";
						WHEN "0000001010111000" =>
						DD(7, 20) <= packet_in;
						counter <= "0000001010111001";
						WHEN "0000001010111001" =>
						DD(7, 21) <= packet_in;
						counter <= "0000001010111010";
						WHEN "0000001010111010" =>
						DD(7, 22) <= packet_in;
						counter <= "0000001010111011";
						WHEN "0000001010111011" =>
						DD(7, 23) <= packet_in;
						counter <= "0000001010111100";
						WHEN "0000001010111100" =>
						DD(7, 24) <= packet_in;
						counter <= "0000001010111101";
						WHEN "0000001010111101" =>
						DD(7, 25) <= packet_in;
						counter <= "0000001010111110";
						WHEN "0000001010111110" =>
						DD(7, 26) <= packet_in;
						counter <= "0000001010111111";
						WHEN "0000001010111111" =>
						DD(7, 27) <= packet_in;
						counter <= "0000001011000000";
						WHEN "0000001011000000" =>
						DD(7, 28) <= packet_in;
						counter <= "0000001011000001";
						WHEN "0000001011000001" =>
						DD(7, 29) <= packet_in;
						counter <= "0000001011000010";
						WHEN "0000001011000010" =>
						DD(7, 30) <= packet_in;
						counter <= "0000001011000011";
						WHEN "0000001011000011" =>
						DD(7, 31) <= packet_in;
						counter <= "0000001011000100";
						WHEN "0000001011000100" =>
						DD(7, 32) <= packet_in;
						counter <= "0000001011000101";
						WHEN "0000001011000101" =>
						DD(7, 33) <= packet_in;
						counter <= "0000001011000110";
						WHEN "0000001011000110" =>
						DD(7, 34) <= packet_in;
						counter <= "0000001011000111";
						WHEN "0000001011000111" =>
						DD(7, 35) <= packet_in;
						counter <= "0000001011001000";
						WHEN "0000001011001000" =>
						DD(7, 36) <= packet_in;
						counter <= "0000001011001001";
						WHEN "0000001011001001" =>
						DD(7, 37) <= packet_in;
						counter <= "0000001011001010";
						WHEN "0000001011001010" =>
						DD(7, 38) <= packet_in;
						counter <= "0000001011001011";
						WHEN "0000001011001011" =>
						DD(7, 39) <= packet_in;
						counter <= "0000001011001100";
						WHEN "0000001011001100" =>
						DD(7, 40) <= packet_in;
						counter <= "0000001011001101";
						WHEN "0000001011001101" =>
						DD(7, 41) <= packet_in;
						counter <= "0000001011001110";
						WHEN "0000001011001110" =>
						DD(7, 42) <= packet_in;
						counter <= "0000001011001111";
						WHEN "0000001011001111" =>
						DD(7, 43) <= packet_in;
						counter <= "0000001011010000";
						WHEN "0000001011010000" =>
						DD(7, 44) <= packet_in;
						counter <= "0000001011010001";
						WHEN "0000001011010001" =>
						DD(7, 45) <= packet_in;
						counter <= "0000001011010010";
						WHEN "0000001011010010" =>
						DD(7, 46) <= packet_in;
						counter <= "0000001011010011";
						WHEN "0000001011010011" =>
						DD(7, 47) <= packet_in;
						counter <= "0000001011010100";
						WHEN "0000001011010100" =>
						DD(7, 48) <= packet_in;
						counter <= "0000001011010101";
						WHEN "0000001011010101" =>
						DD(7, 49) <= packet_in;
						counter <= "0000001011010110";
						WHEN "0000001011010110" =>
						DD(7, 50) <= packet_in;
						counter <= "0000001011010111";
						WHEN "0000001011010111" =>
						DD(7, 51) <= packet_in;
						counter <= "0000001011011000";
						WHEN "0000001011011000" =>
						DD(7, 52) <= packet_in;
						counter <= "0000001011011001";
						WHEN "0000001011011001" =>
						DD(7, 53) <= packet_in;
						counter <= "0000001011011010";
						WHEN "0000001011011010" =>
						DD(7, 54) <= packet_in;
						counter <= "0000001011011011";
						WHEN "0000001011011011" =>
						DD(7, 55) <= packet_in;
						counter <= "0000001011011100";
						WHEN "0000001011011100" =>
						DD(7, 56) <= packet_in;
						counter <= "0000001011011101";
						WHEN "0000001011011101" =>
						DD(7, 57) <= packet_in;
						counter <= "0000001011011110";
						WHEN "0000001011011110" =>
						DD(7, 58) <= packet_in;
						counter <= "0000001011011111";
						WHEN "0000001011011111" =>
						DD(7, 59) <= packet_in;
						counter <= "0000001011100000";
						WHEN "0000001011100000" =>
						DD(7, 60) <= packet_in;
						counter <= "0000001011100001";
						WHEN "0000001011100001" =>
						DD(7, 61) <= packet_in;
						counter <= "0000001011100010";
						WHEN "0000001011100010" =>
						DD(7, 62) <= packet_in;
						counter <= "0000001011100011";
						WHEN "0000001011100011" =>
						DD(7, 63) <= packet_in;
						counter <= "0000001011100100";
						WHEN "0000001011100100" =>
						DD(7, 64) <= packet_in;
						counter <= "0000001011100101";
						WHEN "0000001011100101" =>
						DD(7, 65) <= packet_in;
						counter <= "0000001011100110";
						WHEN "0000001011100110" =>
						DD(7, 66) <= packet_in;
						counter <= "0000001011100111";
						WHEN "0000001011100111" =>
						DD(7, 67) <= packet_in;
						counter <= "0000001011101000";
						WHEN "0000001011101000" =>
						DD(7, 68) <= packet_in;
						counter <= "0000001011101001";
						WHEN "0000001011101001" =>
						DD(7, 69) <= packet_in;
						counter <= "0000001011101010";
						WHEN "0000001011101010" =>
						DD(7, 70) <= packet_in;
						counter <= "0000001011101011";
						WHEN "0000001011101011" =>
						DD(7, 71) <= packet_in;
						counter <= "0000001011101100";
						WHEN "0000001011101100" =>
						DD(7, 72) <= packet_in;
						counter <= "0000001011101101";
						WHEN "0000001011101101" =>
						DD(7, 73) <= packet_in;
						counter <= "0000001011101110";
						WHEN "0000001011101110" =>
						DD(7, 74) <= packet_in;
						counter <= "0000001011101111";
						WHEN "0000001011101111" =>
						DD(7, 75) <= packet_in;
						counter <= "0000001011110000";
						WHEN "0000001011110000" =>
						DD(7, 76) <= packet_in;
						counter <= "0000001011110001";
						WHEN "0000001011110001" =>
						DD(7, 77) <= packet_in;
						counter <= "0000001011110010";
						WHEN "0000001011110010" =>
						DD(7, 78) <= packet_in;
						counter <= "0000001011110011";
						WHEN "0000001011110011" =>
						DD(7, 79) <= packet_in;
						counter <= "0000001011110100";
						WHEN "0000001011110100" =>
						DD(7, 80) <= packet_in;
						counter <= "0000001011110101";
						WHEN "0000001011110101" =>
						DD(7, 81) <= packet_in;
						counter <= "0000001011110110";
						WHEN "0000001011110110" =>
						DD(7, 82) <= packet_in;
						counter <= "0000001011110111";
						WHEN "0000001011110111" =>
						DD(7, 83) <= packet_in;
						counter <= "0000001011111000";
						WHEN "0000001011111000" =>
						DD(7, 84) <= packet_in;
						counter <= "0000001011111001";
						WHEN "0000001011111001" =>
						DD(7, 85) <= packet_in;
						counter <= "0000001011111010";
						WHEN "0000001011111010" =>
						DD(7, 86) <= packet_in;
						counter <= "0000001011111011";
						WHEN "0000001011111011" =>
						DD(7, 87) <= packet_in;
						counter <= "0000001011111100";
						WHEN "0000001011111100" =>
						DD(7, 88) <= packet_in;
						counter <= "0000001011111101";
						WHEN "0000001011111101" =>
						DD(7, 89) <= packet_in;
						counter <= "0000001011111110";
						WHEN "0000001011111110" =>
						DD(7, 90) <= packet_in;
						counter <= "0000001011111111";
						WHEN "0000001011111111" =>
						DD(7, 91) <= packet_in;
						counter <= "0000001100000000";
						WHEN "0000001100000000" =>
						DD(8, 0) <= packet_in;
						counter <= "0000001100000001";
						WHEN "0000001100000001" =>
						DD(8, 1) <= packet_in;
						counter <= "0000001100000010";
						WHEN "0000001100000010" =>
						DD(8, 2) <= packet_in;
						counter <= "0000001100000011";
						WHEN "0000001100000011" =>
						DD(8, 3) <= packet_in;
						counter <= "0000001100000100";
						WHEN "0000001100000100" =>
						DD(8, 4) <= packet_in;
						counter <= "0000001100000101";
						WHEN "0000001100000101" =>
						DD(8, 5) <= packet_in;
						counter <= "0000001100000110";
						WHEN "0000001100000110" =>
						DD(8, 6) <= packet_in;
						counter <= "0000001100000111";
						WHEN "0000001100000111" =>
						DD(8, 7) <= packet_in;
						counter <= "0000001100001000";
						WHEN "0000001100001000" =>
						DD(8, 8) <= packet_in;
						counter <= "0000001100001001";
						WHEN "0000001100001001" =>
						DD(8, 9) <= packet_in;
						counter <= "0000001100001010";
						WHEN "0000001100001010" =>
						DD(8, 10) <= packet_in;
						counter <= "0000001100001011";
						WHEN "0000001100001011" =>
						DD(8, 11) <= packet_in;
						counter <= "0000001100001100";
						WHEN "0000001100001100" =>
						DD(8, 12) <= packet_in;
						counter <= "0000001100001101";
						WHEN "0000001100001101" =>
						DD(8, 13) <= packet_in;
						counter <= "0000001100001110";
						WHEN "0000001100001110" =>
						DD(8, 14) <= packet_in;
						counter <= "0000001100001111";
						WHEN "0000001100001111" =>
						DD(8, 15) <= packet_in;
						counter <= "0000001100010000";
						WHEN "0000001100010000" =>
						DD(8, 16) <= packet_in;
						counter <= "0000001100010001";
						WHEN "0000001100010001" =>
						DD(8, 17) <= packet_in;
						counter <= "0000001100010010";
						WHEN "0000001100010010" =>
						DD(8, 18) <= packet_in;
						counter <= "0000001100010011";
						WHEN "0000001100010011" =>
						DD(8, 19) <= packet_in;
						counter <= "0000001100010100";
						WHEN "0000001100010100" =>
						DD(8, 20) <= packet_in;
						counter <= "0000001100010101";
						WHEN "0000001100010101" =>
						DD(8, 21) <= packet_in;
						counter <= "0000001100010110";
						WHEN "0000001100010110" =>
						DD(8, 22) <= packet_in;
						counter <= "0000001100010111";
						WHEN "0000001100010111" =>
						DD(8, 23) <= packet_in;
						counter <= "0000001100011000";
						WHEN "0000001100011000" =>
						DD(8, 24) <= packet_in;
						counter <= "0000001100011001";
						WHEN "0000001100011001" =>
						DD(8, 25) <= packet_in;
						counter <= "0000001100011010";
						WHEN "0000001100011010" =>
						DD(8, 26) <= packet_in;
						counter <= "0000001100011011";
						WHEN "0000001100011011" =>
						DD(8, 27) <= packet_in;
						counter <= "0000001100011100";
						WHEN "0000001100011100" =>
						DD(8, 28) <= packet_in;
						counter <= "0000001100011101";
						WHEN "0000001100011101" =>
						DD(8, 29) <= packet_in;
						counter <= "0000001100011110";
						WHEN "0000001100011110" =>
						DD(8, 30) <= packet_in;
						counter <= "0000001100011111";
						WHEN "0000001100011111" =>
						DD(8, 31) <= packet_in;
						counter <= "0000001100100000";
						WHEN "0000001100100000" =>
						DD(8, 32) <= packet_in;
						counter <= "0000001100100001";
						WHEN "0000001100100001" =>
						DD(8, 33) <= packet_in;
						counter <= "0000001100100010";
						WHEN "0000001100100010" =>
						DD(8, 34) <= packet_in;
						counter <= "0000001100100011";
						WHEN "0000001100100011" =>
						DD(8, 35) <= packet_in;
						counter <= "0000001100100100";
						WHEN "0000001100100100" =>
						DD(8, 36) <= packet_in;
						counter <= "0000001100100101";
						WHEN "0000001100100101" =>
						DD(8, 37) <= packet_in;
						counter <= "0000001100100110";
						WHEN "0000001100100110" =>
						DD(8, 38) <= packet_in;
						counter <= "0000001100100111";
						WHEN "0000001100100111" =>
						DD(8, 39) <= packet_in;
						counter <= "0000001100101000";
						WHEN "0000001100101000" =>
						DD(8, 40) <= packet_in;
						counter <= "0000001100101001";
						WHEN "0000001100101001" =>
						DD(8, 41) <= packet_in;
						counter <= "0000001100101010";
						WHEN "0000001100101010" =>
						DD(8, 42) <= packet_in;
						counter <= "0000001100101011";
						WHEN "0000001100101011" =>
						DD(8, 43) <= packet_in;
						counter <= "0000001100101100";
						WHEN "0000001100101100" =>
						DD(8, 44) <= packet_in;
						counter <= "0000001100101101";
						WHEN "0000001100101101" =>
						DD(8, 45) <= packet_in;
						counter <= "0000001100101110";
						WHEN "0000001100101110" =>
						DD(8, 46) <= packet_in;
						counter <= "0000001100101111";
						WHEN "0000001100101111" =>
						DD(8, 47) <= packet_in;
						counter <= "0000001100110000";
						WHEN "0000001100110000" =>
						DD(8, 48) <= packet_in;
						counter <= "0000001100110001";
						WHEN "0000001100110001" =>
						DD(8, 49) <= packet_in;
						counter <= "0000001100110010";
						WHEN "0000001100110010" =>
						DD(8, 50) <= packet_in;
						counter <= "0000001100110011";
						WHEN "0000001100110011" =>
						DD(8, 51) <= packet_in;
						counter <= "0000001100110100";
						WHEN "0000001100110100" =>
						DD(8, 52) <= packet_in;
						counter <= "0000001100110101";
						WHEN "0000001100110101" =>
						DD(8, 53) <= packet_in;
						counter <= "0000001100110110";
						WHEN "0000001100110110" =>
						DD(8, 54) <= packet_in;
						counter <= "0000001100110111";
						WHEN "0000001100110111" =>
						DD(8, 55) <= packet_in;
						counter <= "0000001100111000";
						WHEN "0000001100111000" =>
						DD(8, 56) <= packet_in;
						counter <= "0000001100111001";
						WHEN "0000001100111001" =>
						DD(8, 57) <= packet_in;
						counter <= "0000001100111010";
						WHEN "0000001100111010" =>
						DD(8, 58) <= packet_in;
						counter <= "0000001100111011";
						WHEN "0000001100111011" =>
						DD(8, 59) <= packet_in;
						counter <= "0000001100111100";
						WHEN "0000001100111100" =>
						DD(8, 60) <= packet_in;
						counter <= "0000001100111101";
						WHEN "0000001100111101" =>
						DD(8, 61) <= packet_in;
						counter <= "0000001100111110";
						WHEN "0000001100111110" =>
						DD(8, 62) <= packet_in;
						counter <= "0000001100111111";
						WHEN "0000001100111111" =>
						DD(8, 63) <= packet_in;
						counter <= "0000001101000000";
						WHEN "0000001101000000" =>
						DD(8, 64) <= packet_in;
						counter <= "0000001101000001";
						WHEN "0000001101000001" =>
						DD(8, 65) <= packet_in;
						counter <= "0000001101000010";
						WHEN "0000001101000010" =>
						DD(8, 66) <= packet_in;
						counter <= "0000001101000011";
						WHEN "0000001101000011" =>
						DD(8, 67) <= packet_in;
						counter <= "0000001101000100";
						WHEN "0000001101000100" =>
						DD(8, 68) <= packet_in;
						counter <= "0000001101000101";
						WHEN "0000001101000101" =>
						DD(8, 69) <= packet_in;
						counter <= "0000001101000110";
						WHEN "0000001101000110" =>
						DD(8, 70) <= packet_in;
						counter <= "0000001101000111";
						WHEN "0000001101000111" =>
						DD(8, 71) <= packet_in;
						counter <= "0000001101001000";
						WHEN "0000001101001000" =>
						DD(8, 72) <= packet_in;
						counter <= "0000001101001001";
						WHEN "0000001101001001" =>
						DD(8, 73) <= packet_in;
						counter <= "0000001101001010";
						WHEN "0000001101001010" =>
						DD(8, 74) <= packet_in;
						counter <= "0000001101001011";
						WHEN "0000001101001011" =>
						DD(8, 75) <= packet_in;
						counter <= "0000001101001100";
						WHEN "0000001101001100" =>
						DD(8, 76) <= packet_in;
						counter <= "0000001101001101";
						WHEN "0000001101001101" =>
						DD(8, 77) <= packet_in;
						counter <= "0000001101001110";
						WHEN "0000001101001110" =>
						DD(8, 78) <= packet_in;
						counter <= "0000001101001111";
						WHEN "0000001101001111" =>
						DD(8, 79) <= packet_in;
						counter <= "0000001101010000";
						WHEN "0000001101010000" =>
						DD(8, 80) <= packet_in;
						counter <= "0000001101010001";
						WHEN "0000001101010001" =>
						DD(8, 81) <= packet_in;
						counter <= "0000001101010010";
						WHEN "0000001101010010" =>
						DD(8, 82) <= packet_in;
						counter <= "0000001101010011";
						WHEN "0000001101010011" =>
						DD(8, 83) <= packet_in;
						counter <= "0000001101010100";
						WHEN "0000001101010100" =>
						DD(8, 84) <= packet_in;
						counter <= "0000001101010101";
						WHEN "0000001101010101" =>
						DD(8, 85) <= packet_in;
						counter <= "0000001101010110";
						WHEN "0000001101010110" =>
						DD(8, 86) <= packet_in;
						counter <= "0000001101010111";
						WHEN "0000001101010111" =>
						DD(8, 87) <= packet_in;
						counter <= "0000001101011000";
						WHEN "0000001101011000" =>
						DD(8, 88) <= packet_in;
						counter <= "0000001101011001";
						WHEN "0000001101011001" =>
						DD(8, 89) <= packet_in;
						counter <= "0000001101011010";
						WHEN "0000001101011010" =>
						DD(8, 90) <= packet_in;
						counter <= "0000001101011011";
						WHEN "0000001101011011" =>
						DD(8, 91) <= packet_in;
						counter <= "0000001101011100";
						WHEN "0000001101011100" =>
						DD(9, 0) <= packet_in;
						counter <= "0000001101011101";
						WHEN "0000001101011101" =>
						DD(9, 1) <= packet_in;
						counter <= "0000001101011110";
						WHEN "0000001101011110" =>
						DD(9, 2) <= packet_in;
						counter <= "0000001101011111";
						WHEN "0000001101011111" =>
						DD(9, 3) <= packet_in;
						counter <= "0000001101100000";
						WHEN "0000001101100000" =>
						DD(9, 4) <= packet_in;
						counter <= "0000001101100001";
						WHEN "0000001101100001" =>
						DD(9, 5) <= packet_in;
						counter <= "0000001101100010";
						WHEN "0000001101100010" =>
						DD(9, 6) <= packet_in;
						counter <= "0000001101100011";
						WHEN "0000001101100011" =>
						DD(9, 7) <= packet_in;
						counter <= "0000001101100100";
						WHEN "0000001101100100" =>
						DD(9, 8) <= packet_in;
						counter <= "0000001101100101";
						WHEN "0000001101100101" =>
						DD(9, 9) <= packet_in;
						counter <= "0000001101100110";
						WHEN "0000001101100110" =>
						DD(9, 10) <= packet_in;
						counter <= "0000001101100111";
						WHEN "0000001101100111" =>
						DD(9, 11) <= packet_in;
						counter <= "0000001101101000";
						WHEN "0000001101101000" =>
						DD(9, 12) <= packet_in;
						counter <= "0000001101101001";
						WHEN "0000001101101001" =>
						DD(9, 13) <= packet_in;
						counter <= "0000001101101010";
						WHEN "0000001101101010" =>
						DD(9, 14) <= packet_in;
						counter <= "0000001101101011";
						WHEN "0000001101101011" =>
						DD(9, 15) <= packet_in;
						counter <= "0000001101101100";
						WHEN "0000001101101100" =>
						DD(9, 16) <= packet_in;
						counter <= "0000001101101101";
						WHEN "0000001101101101" =>
						DD(9, 17) <= packet_in;
						counter <= "0000001101101110";
						WHEN "0000001101101110" =>
						DD(9, 18) <= packet_in;
						counter <= "0000001101101111";
						WHEN "0000001101101111" =>
						DD(9, 19) <= packet_in;
						counter <= "0000001101110000";
						WHEN "0000001101110000" =>
						DD(9, 20) <= packet_in;
						counter <= "0000001101110001";
						WHEN "0000001101110001" =>
						DD(9, 21) <= packet_in;
						counter <= "0000001101110010";
						WHEN "0000001101110010" =>
						DD(9, 22) <= packet_in;
						counter <= "0000001101110011";
						WHEN "0000001101110011" =>
						DD(9, 23) <= packet_in;
						counter <= "0000001101110100";
						WHEN "0000001101110100" =>
						DD(9, 24) <= packet_in;
						counter <= "0000001101110101";
						WHEN "0000001101110101" =>
						DD(9, 25) <= packet_in;
						counter <= "0000001101110110";
						WHEN "0000001101110110" =>
						DD(9, 26) <= packet_in;
						counter <= "0000001101110111";
						WHEN "0000001101110111" =>
						DD(9, 27) <= packet_in;
						counter <= "0000001101111000";
						WHEN "0000001101111000" =>
						DD(9, 28) <= packet_in;
						counter <= "0000001101111001";
						WHEN "0000001101111001" =>
						DD(9, 29) <= packet_in;
						counter <= "0000001101111010";
						WHEN "0000001101111010" =>
						DD(9, 30) <= packet_in;
						counter <= "0000001101111011";
						WHEN "0000001101111011" =>
						DD(9, 31) <= packet_in;
						counter <= "0000001101111100";
						WHEN "0000001101111100" =>
						DD(9, 32) <= packet_in;
						counter <= "0000001101111101";
						WHEN "0000001101111101" =>
						DD(9, 33) <= packet_in;
						counter <= "0000001101111110";
						WHEN "0000001101111110" =>
						DD(9, 34) <= packet_in;
						counter <= "0000001101111111";
						WHEN "0000001101111111" =>
						DD(9, 35) <= packet_in;
						counter <= "0000001110000000";
						WHEN "0000001110000000" =>
						DD(9, 36) <= packet_in;
						counter <= "0000001110000001";
						WHEN "0000001110000001" =>
						DD(9, 37) <= packet_in;
						counter <= "0000001110000010";
						WHEN "0000001110000010" =>
						DD(9, 38) <= packet_in;
						counter <= "0000001110000011";
						WHEN "0000001110000011" =>
						DD(9, 39) <= packet_in;
						counter <= "0000001110000100";
						WHEN "0000001110000100" =>
						DD(9, 40) <= packet_in;
						counter <= "0000001110000101";
						WHEN "0000001110000101" =>
						DD(9, 41) <= packet_in;
						counter <= "0000001110000110";
						WHEN "0000001110000110" =>
						DD(9, 42) <= packet_in;
						counter <= "0000001110000111";
						WHEN "0000001110000111" =>
						DD(9, 43) <= packet_in;
						counter <= "0000001110001000";
						WHEN "0000001110001000" =>
						DD(9, 44) <= packet_in;
						counter <= "0000001110001001";
						WHEN "0000001110001001" =>
						DD(9, 45) <= packet_in;
						counter <= "0000001110001010";
						WHEN "0000001110001010" =>
						DD(9, 46) <= packet_in;
						counter <= "0000001110001011";
						WHEN "0000001110001011" =>
						DD(9, 47) <= packet_in;
						counter <= "0000001110001100";
						WHEN "0000001110001100" =>
						DD(9, 48) <= packet_in;
						counter <= "0000001110001101";
						WHEN "0000001110001101" =>
						DD(9, 49) <= packet_in;
						counter <= "0000001110001110";
						WHEN "0000001110001110" =>
						DD(9, 50) <= packet_in;
						counter <= "0000001110001111";
						WHEN "0000001110001111" =>
						DD(9, 51) <= packet_in;
						counter <= "0000001110010000";
						WHEN "0000001110010000" =>
						DD(9, 52) <= packet_in;
						counter <= "0000001110010001";
						WHEN "0000001110010001" =>
						DD(9, 53) <= packet_in;
						counter <= "0000001110010010";
						WHEN "0000001110010010" =>
						DD(9, 54) <= packet_in;
						counter <= "0000001110010011";
						WHEN "0000001110010011" =>
						DD(9, 55) <= packet_in;
						counter <= "0000001110010100";
						WHEN "0000001110010100" =>
						DD(9, 56) <= packet_in;
						counter <= "0000001110010101";
						WHEN "0000001110010101" =>
						DD(9, 57) <= packet_in;
						counter <= "0000001110010110";
						WHEN "0000001110010110" =>
						DD(9, 58) <= packet_in;
						counter <= "0000001110010111";
						WHEN "0000001110010111" =>
						DD(9, 59) <= packet_in;
						counter <= "0000001110011000";
						WHEN "0000001110011000" =>
						DD(9, 60) <= packet_in;
						counter <= "0000001110011001";
						WHEN "0000001110011001" =>
						DD(9, 61) <= packet_in;
						counter <= "0000001110011010";
						WHEN "0000001110011010" =>
						DD(9, 62) <= packet_in;
						counter <= "0000001110011011";
						WHEN "0000001110011011" =>
						DD(9, 63) <= packet_in;
						counter <= "0000001110011100";
						WHEN "0000001110011100" =>
						DD(9, 64) <= packet_in;
						counter <= "0000001110011101";
						WHEN "0000001110011101" =>
						DD(9, 65) <= packet_in;
						counter <= "0000001110011110";
						WHEN "0000001110011110" =>
						DD(9, 66) <= packet_in;
						counter <= "0000001110011111";
						WHEN "0000001110011111" =>
						DD(9, 67) <= packet_in;
						counter <= "0000001110100000";
						WHEN "0000001110100000" =>
						DD(9, 68) <= packet_in;
						counter <= "0000001110100001";
						WHEN "0000001110100001" =>
						DD(9, 69) <= packet_in;
						counter <= "0000001110100010";
						WHEN "0000001110100010" =>
						DD(9, 70) <= packet_in;
						counter <= "0000001110100011";
						WHEN "0000001110100011" =>
						DD(9, 71) <= packet_in;
						counter <= "0000001110100100";
						WHEN "0000001110100100" =>
						DD(9, 72) <= packet_in;
						counter <= "0000001110100101";
						WHEN "0000001110100101" =>
						DD(9, 73) <= packet_in;
						counter <= "0000001110100110";
						WHEN "0000001110100110" =>
						DD(9, 74) <= packet_in;
						counter <= "0000001110100111";
						WHEN "0000001110100111" =>
						DD(9, 75) <= packet_in;
						counter <= "0000001110101000";
						WHEN "0000001110101000" =>
						DD(9, 76) <= packet_in;
						counter <= "0000001110101001";
						WHEN "0000001110101001" =>
						DD(9, 77) <= packet_in;
						counter <= "0000001110101010";
						WHEN "0000001110101010" =>
						DD(9, 78) <= packet_in;
						counter <= "0000001110101011";
						WHEN "0000001110101011" =>
						DD(9, 79) <= packet_in;
						counter <= "0000001110101100";
						WHEN "0000001110101100" =>
						DD(9, 80) <= packet_in;
						counter <= "0000001110101101";
						WHEN "0000001110101101" =>
						DD(9, 81) <= packet_in;
						counter <= "0000001110101110";
						WHEN "0000001110101110" =>
						DD(9, 82) <= packet_in;
						counter <= "0000001110101111";
						WHEN "0000001110101111" =>
						DD(9, 83) <= packet_in;
						counter <= "0000001110110000";
						WHEN "0000001110110000" =>
						DD(9, 84) <= packet_in;
						counter <= "0000001110110001";
						WHEN "0000001110110001" =>
						DD(9, 85) <= packet_in;
						counter <= "0000001110110010";
						WHEN "0000001110110010" =>
						DD(9, 86) <= packet_in;
						counter <= "0000001110110011";
						WHEN "0000001110110011" =>
						DD(9, 87) <= packet_in;
						counter <= "0000001110110100";
						WHEN "0000001110110100" =>
						DD(9, 88) <= packet_in;
						counter <= "0000001110110101";
						WHEN "0000001110110101" =>
						DD(9, 89) <= packet_in;
						counter <= "0000001110110110";
						WHEN "0000001110110110" =>
						DD(9, 90) <= packet_in;
						counter <= "0000001110110111";
						WHEN "0000001110110111" =>
						DD(9, 91) <= packet_in;
						counter <= "0000001110111000";
						WHEN "0000001110111000" =>
						DD(10, 0) <= packet_in;
						counter <= "0000001110111001";
						WHEN "0000001110111001" =>
						DD(10, 1) <= packet_in;
						counter <= "0000001110111010";
						WHEN "0000001110111010" =>
						DD(10, 2) <= packet_in;
						counter <= "0000001110111011";
						WHEN "0000001110111011" =>
						DD(10, 3) <= packet_in;
						counter <= "0000001110111100";
						WHEN "0000001110111100" =>
						DD(10, 4) <= packet_in;
						counter <= "0000001110111101";
						WHEN "0000001110111101" =>
						DD(10, 5) <= packet_in;
						counter <= "0000001110111110";
						WHEN "0000001110111110" =>
						DD(10, 6) <= packet_in;
						counter <= "0000001110111111";
						WHEN "0000001110111111" =>
						DD(10, 7) <= packet_in;
						counter <= "0000001111000000";
						WHEN "0000001111000000" =>
						DD(10, 8) <= packet_in;
						counter <= "0000001111000001";
						WHEN "0000001111000001" =>
						DD(10, 9) <= packet_in;
						counter <= "0000001111000010";
						WHEN "0000001111000010" =>
						DD(10, 10) <= packet_in;
						counter <= "0000001111000011";
						WHEN "0000001111000011" =>
						DD(10, 11) <= packet_in;
						counter <= "0000001111000100";
						WHEN "0000001111000100" =>
						DD(10, 12) <= packet_in;
						counter <= "0000001111000101";
						WHEN "0000001111000101" =>
						DD(10, 13) <= packet_in;
						counter <= "0000001111000110";
						WHEN "0000001111000110" =>
						DD(10, 14) <= packet_in;
						counter <= "0000001111000111";
						WHEN "0000001111000111" =>
						DD(10, 15) <= packet_in;
						counter <= "0000001111001000";
						WHEN "0000001111001000" =>
						DD(10, 16) <= packet_in;
						counter <= "0000001111001001";
						WHEN "0000001111001001" =>
						DD(10, 17) <= packet_in;
						counter <= "0000001111001010";
						WHEN "0000001111001010" =>
						DD(10, 18) <= packet_in;
						counter <= "0000001111001011";
						WHEN "0000001111001011" =>
						DD(10, 19) <= packet_in;
						counter <= "0000001111001100";
						WHEN "0000001111001100" =>
						DD(10, 20) <= packet_in;
						counter <= "0000001111001101";
						WHEN "0000001111001101" =>
						DD(10, 21) <= packet_in;
						counter <= "0000001111001110";
						WHEN "0000001111001110" =>
						DD(10, 22) <= packet_in;
						counter <= "0000001111001111";
						WHEN "0000001111001111" =>
						DD(10, 23) <= packet_in;
						counter <= "0000001111010000";
						WHEN "0000001111010000" =>
						DD(10, 24) <= packet_in;
						counter <= "0000001111010001";
						WHEN "0000001111010001" =>
						DD(10, 25) <= packet_in;
						counter <= "0000001111010010";
						WHEN "0000001111010010" =>
						DD(10, 26) <= packet_in;
						counter <= "0000001111010011";
						WHEN "0000001111010011" =>
						DD(10, 27) <= packet_in;
						counter <= "0000001111010100";
						WHEN "0000001111010100" =>
						DD(10, 28) <= packet_in;
						counter <= "0000001111010101";
						WHEN "0000001111010101" =>
						DD(10, 29) <= packet_in;
						counter <= "0000001111010110";
						WHEN "0000001111010110" =>
						DD(10, 30) <= packet_in;
						counter <= "0000001111010111";
						WHEN "0000001111010111" =>
						DD(10, 31) <= packet_in;
						counter <= "0000001111011000";
						WHEN "0000001111011000" =>
						DD(10, 32) <= packet_in;
						counter <= "0000001111011001";
						WHEN "0000001111011001" =>
						DD(10, 33) <= packet_in;
						counter <= "0000001111011010";
						WHEN "0000001111011010" =>
						DD(10, 34) <= packet_in;
						counter <= "0000001111011011";
						WHEN "0000001111011011" =>
						DD(10, 35) <= packet_in;
						counter <= "0000001111011100";
						WHEN "0000001111011100" =>
						DD(10, 36) <= packet_in;
						counter <= "0000001111011101";
						WHEN "0000001111011101" =>
						DD(10, 37) <= packet_in;
						counter <= "0000001111011110";
						WHEN "0000001111011110" =>
						DD(10, 38) <= packet_in;
						counter <= "0000001111011111";
						WHEN "0000001111011111" =>
						DD(10, 39) <= packet_in;
						counter <= "0000001111100000";
						WHEN "0000001111100000" =>
						DD(10, 40) <= packet_in;
						counter <= "0000001111100001";
						WHEN "0000001111100001" =>
						DD(10, 41) <= packet_in;
						counter <= "0000001111100010";
						WHEN "0000001111100010" =>
						DD(10, 42) <= packet_in;
						counter <= "0000001111100011";
						WHEN "0000001111100011" =>
						DD(10, 43) <= packet_in;
						counter <= "0000001111100100";
						WHEN "0000001111100100" =>
						DD(10, 44) <= packet_in;
						counter <= "0000001111100101";
						WHEN "0000001111100101" =>
						DD(10, 45) <= packet_in;
						counter <= "0000001111100110";
						WHEN "0000001111100110" =>
						DD(10, 46) <= packet_in;
						counter <= "0000001111100111";
						WHEN "0000001111100111" =>
						DD(10, 47) <= packet_in;
						counter <= "0000001111101000";
						WHEN "0000001111101000" =>
						DD(10, 48) <= packet_in;
						counter <= "0000001111101001";
						WHEN "0000001111101001" =>
						DD(10, 49) <= packet_in;
						counter <= "0000001111101010";
						WHEN "0000001111101010" =>
						DD(10, 50) <= packet_in;
						counter <= "0000001111101011";
						WHEN "0000001111101011" =>
						DD(10, 51) <= packet_in;
						counter <= "0000001111101100";
						WHEN "0000001111101100" =>
						DD(10, 52) <= packet_in;
						counter <= "0000001111101101";
						WHEN "0000001111101101" =>
						DD(10, 53) <= packet_in;
						counter <= "0000001111101110";
						WHEN "0000001111101110" =>
						DD(10, 54) <= packet_in;
						counter <= "0000001111101111";
						WHEN "0000001111101111" =>
						DD(10, 55) <= packet_in;
						counter <= "0000001111110000";
						WHEN "0000001111110000" =>
						DD(10, 56) <= packet_in;
						counter <= "0000001111110001";
						WHEN "0000001111110001" =>
						DD(10, 57) <= packet_in;
						counter <= "0000001111110010";
						WHEN "0000001111110010" =>
						DD(10, 58) <= packet_in;
						counter <= "0000001111110011";
						WHEN "0000001111110011" =>
						DD(10, 59) <= packet_in;
						counter <= "0000001111110100";
						WHEN "0000001111110100" =>
						DD(10, 60) <= packet_in;
						counter <= "0000001111110101";
						WHEN "0000001111110101" =>
						DD(10, 61) <= packet_in;
						counter <= "0000001111110110";
						WHEN "0000001111110110" =>
						DD(10, 62) <= packet_in;
						counter <= "0000001111110111";
						WHEN "0000001111110111" =>
						DD(10, 63) <= packet_in;
						counter <= "0000001111111000";
						WHEN "0000001111111000" =>
						DD(10, 64) <= packet_in;
						counter <= "0000001111111001";
						WHEN "0000001111111001" =>
						DD(10, 65) <= packet_in;
						counter <= "0000001111111010";
						WHEN "0000001111111010" =>
						DD(10, 66) <= packet_in;
						counter <= "0000001111111011";
						WHEN "0000001111111011" =>
						DD(10, 67) <= packet_in;
						counter <= "0000001111111100";
						WHEN "0000001111111100" =>
						DD(10, 68) <= packet_in;
						counter <= "0000001111111101";
						WHEN "0000001111111101" =>
						DD(10, 69) <= packet_in;
						counter <= "0000001111111110";
						WHEN "0000001111111110" =>
						DD(10, 70) <= packet_in;
						counter <= "0000001111111111";
						WHEN "0000001111111111" =>
						DD(10, 71) <= packet_in;
						counter <= "0000010000000000";
						WHEN "0000010000000000" =>
						DD(10, 72) <= packet_in;
						counter <= "0000010000000001";
						WHEN "0000010000000001" =>
						DD(10, 73) <= packet_in;
						counter <= "0000010000000010";
						WHEN "0000010000000010" =>
						DD(10, 74) <= packet_in;
						counter <= "0000010000000011";
						WHEN "0000010000000011" =>
						DD(10, 75) <= packet_in;
						counter <= "0000010000000100";
						WHEN "0000010000000100" =>
						DD(10, 76) <= packet_in;
						counter <= "0000010000000101";
						WHEN "0000010000000101" =>
						DD(10, 77) <= packet_in;
						counter <= "0000010000000110";
						WHEN "0000010000000110" =>
						DD(10, 78) <= packet_in;
						counter <= "0000010000000111";
						WHEN "0000010000000111" =>
						DD(10, 79) <= packet_in;
						counter <= "0000010000001000";
						WHEN "0000010000001000" =>
						DD(10, 80) <= packet_in;
						counter <= "0000010000001001";
						WHEN "0000010000001001" =>
						DD(10, 81) <= packet_in;
						counter <= "0000010000001010";
						WHEN "0000010000001010" =>
						DD(10, 82) <= packet_in;
						counter <= "0000010000001011";
						WHEN "0000010000001011" =>
						DD(10, 83) <= packet_in;
						counter <= "0000010000001100";
						WHEN "0000010000001100" =>
						DD(10, 84) <= packet_in;
						counter <= "0000010000001101";
						WHEN "0000010000001101" =>
						DD(10, 85) <= packet_in;
						counter <= "0000010000001110";
						WHEN "0000010000001110" =>
						DD(10, 86) <= packet_in;
						counter <= "0000010000001111";
						WHEN "0000010000001111" =>
						DD(10, 87) <= packet_in;
						counter <= "0000010000010000";
						WHEN "0000010000010000" =>
						DD(10, 88) <= packet_in;
						counter <= "0000010000010001";
						WHEN "0000010000010001" =>
						DD(10, 89) <= packet_in;
						counter <= "0000010000010010";
						WHEN "0000010000010010" =>
						DD(10, 90) <= packet_in;
						counter <= "0000010000010011";
						WHEN "0000010000010011" =>
						DD(10, 91) <= packet_in;
						counter <= "0000010000010100";
						WHEN "0000010000010100" =>
						DD(11, 0) <= packet_in;
						counter <= "0000010000010101";
						WHEN "0000010000010101" =>
						DD(11, 1) <= packet_in;
						counter <= "0000010000010110";
						WHEN "0000010000010110" =>
						DD(11, 2) <= packet_in;
						counter <= "0000010000010111";
						WHEN "0000010000010111" =>
						DD(11, 3) <= packet_in;
						counter <= "0000010000011000";
						WHEN "0000010000011000" =>
						DD(11, 4) <= packet_in;
						counter <= "0000010000011001";
						WHEN "0000010000011001" =>
						DD(11, 5) <= packet_in;
						counter <= "0000010000011010";
						WHEN "0000010000011010" =>
						DD(11, 6) <= packet_in;
						counter <= "0000010000011011";
						WHEN "0000010000011011" =>
						DD(11, 7) <= packet_in;
						counter <= "0000010000011100";
						WHEN "0000010000011100" =>
						DD(11, 8) <= packet_in;
						counter <= "0000010000011101";
						WHEN "0000010000011101" =>
						DD(11, 9) <= packet_in;
						counter <= "0000010000011110";
						WHEN "0000010000011110" =>
						DD(11, 10) <= packet_in;
						counter <= "0000010000011111";
						WHEN "0000010000011111" =>
						DD(11, 11) <= packet_in;
						counter <= "0000010000100000";
						WHEN "0000010000100000" =>
						DD(11, 12) <= packet_in;
						counter <= "0000010000100001";
						WHEN "0000010000100001" =>
						DD(11, 13) <= packet_in;
						counter <= "0000010000100010";
						WHEN "0000010000100010" =>
						DD(11, 14) <= packet_in;
						counter <= "0000010000100011";
						WHEN "0000010000100011" =>
						DD(11, 15) <= packet_in;
						counter <= "0000010000100100";
						WHEN "0000010000100100" =>
						DD(11, 16) <= packet_in;
						counter <= "0000010000100101";
						WHEN "0000010000100101" =>
						DD(11, 17) <= packet_in;
						counter <= "0000010000100110";
						WHEN "0000010000100110" =>
						DD(11, 18) <= packet_in;
						counter <= "0000010000100111";
						WHEN "0000010000100111" =>
						DD(11, 19) <= packet_in;
						counter <= "0000010000101000";
						WHEN "0000010000101000" =>
						DD(11, 20) <= packet_in;
						counter <= "0000010000101001";
						WHEN "0000010000101001" =>
						DD(11, 21) <= packet_in;
						counter <= "0000010000101010";
						WHEN "0000010000101010" =>
						DD(11, 22) <= packet_in;
						counter <= "0000010000101011";
						WHEN "0000010000101011" =>
						DD(11, 23) <= packet_in;
						counter <= "0000010000101100";
						WHEN "0000010000101100" =>
						DD(11, 24) <= packet_in;
						counter <= "0000010000101101";
						WHEN "0000010000101101" =>
						DD(11, 25) <= packet_in;
						counter <= "0000010000101110";
						WHEN "0000010000101110" =>
						DD(11, 26) <= packet_in;
						counter <= "0000010000101111";
						WHEN "0000010000101111" =>
						DD(11, 27) <= packet_in;
						counter <= "0000010000110000";
						WHEN "0000010000110000" =>
						DD(11, 28) <= packet_in;
						counter <= "0000010000110001";
						WHEN "0000010000110001" =>
						DD(11, 29) <= packet_in;
						counter <= "0000010000110010";
						WHEN "0000010000110010" =>
						DD(11, 30) <= packet_in;
						counter <= "0000010000110011";
						WHEN "0000010000110011" =>
						DD(11, 31) <= packet_in;
						counter <= "0000010000110100";
						WHEN "0000010000110100" =>
						DD(11, 32) <= packet_in;
						counter <= "0000010000110101";
						WHEN "0000010000110101" =>
						DD(11, 33) <= packet_in;
						counter <= "0000010000110110";
						WHEN "0000010000110110" =>
						DD(11, 34) <= packet_in;
						counter <= "0000010000110111";
						WHEN "0000010000110111" =>
						DD(11, 35) <= packet_in;
						counter <= "0000010000111000";
						WHEN "0000010000111000" =>
						DD(11, 36) <= packet_in;
						counter <= "0000010000111001";
						WHEN "0000010000111001" =>
						DD(11, 37) <= packet_in;
						counter <= "0000010000111010";
						WHEN "0000010000111010" =>
						DD(11, 38) <= packet_in;
						counter <= "0000010000111011";
						WHEN "0000010000111011" =>
						DD(11, 39) <= packet_in;
						counter <= "0000010000111100";
						WHEN "0000010000111100" =>
						DD(11, 40) <= packet_in;
						counter <= "0000010000111101";
						WHEN "0000010000111101" =>
						DD(11, 41) <= packet_in;
						counter <= "0000010000111110";
						WHEN "0000010000111110" =>
						DD(11, 42) <= packet_in;
						counter <= "0000010000111111";
						WHEN "0000010000111111" =>
						DD(11, 43) <= packet_in;
						counter <= "0000010001000000";
						WHEN "0000010001000000" =>
						DD(11, 44) <= packet_in;
						counter <= "0000010001000001";
						WHEN "0000010001000001" =>
						DD(11, 45) <= packet_in;
						counter <= "0000010001000010";
						WHEN "0000010001000010" =>
						DD(11, 46) <= packet_in;
						counter <= "0000010001000011";
						WHEN "0000010001000011" =>
						DD(11, 47) <= packet_in;
						counter <= "0000010001000100";
						WHEN "0000010001000100" =>
						DD(11, 48) <= packet_in;
						counter <= "0000010001000101";
						WHEN "0000010001000101" =>
						DD(11, 49) <= packet_in;
						counter <= "0000010001000110";
						WHEN "0000010001000110" =>
						DD(11, 50) <= packet_in;
						counter <= "0000010001000111";
						WHEN "0000010001000111" =>
						DD(11, 51) <= packet_in;
						counter <= "0000010001001000";
						WHEN "0000010001001000" =>
						DD(11, 52) <= packet_in;
						counter <= "0000010001001001";
						WHEN "0000010001001001" =>
						DD(11, 53) <= packet_in;
						counter <= "0000010001001010";
						WHEN "0000010001001010" =>
						DD(11, 54) <= packet_in;
						counter <= "0000010001001011";
						WHEN "0000010001001011" =>
						DD(11, 55) <= packet_in;
						counter <= "0000010001001100";
						WHEN "0000010001001100" =>
						DD(11, 56) <= packet_in;
						counter <= "0000010001001101";
						WHEN "0000010001001101" =>
						DD(11, 57) <= packet_in;
						counter <= "0000010001001110";
						WHEN "0000010001001110" =>
						DD(11, 58) <= packet_in;
						counter <= "0000010001001111";
						WHEN "0000010001001111" =>
						DD(11, 59) <= packet_in;
						counter <= "0000010001010000";
						WHEN "0000010001010000" =>
						DD(11, 60) <= packet_in;
						counter <= "0000010001010001";
						WHEN "0000010001010001" =>
						DD(11, 61) <= packet_in;
						counter <= "0000010001010010";
						WHEN "0000010001010010" =>
						DD(11, 62) <= packet_in;
						counter <= "0000010001010011";
						WHEN "0000010001010011" =>
						DD(11, 63) <= packet_in;
						counter <= "0000010001010100";
						WHEN "0000010001010100" =>
						DD(11, 64) <= packet_in;
						counter <= "0000010001010101";
						WHEN "0000010001010101" =>
						DD(11, 65) <= packet_in;
						counter <= "0000010001010110";
						WHEN "0000010001010110" =>
						DD(11, 66) <= packet_in;
						counter <= "0000010001010111";
						WHEN "0000010001010111" =>
						DD(11, 67) <= packet_in;
						counter <= "0000010001011000";
						WHEN "0000010001011000" =>
						DD(11, 68) <= packet_in;
						counter <= "0000010001011001";
						WHEN "0000010001011001" =>
						DD(11, 69) <= packet_in;
						counter <= "0000010001011010";
						WHEN "0000010001011010" =>
						DD(11, 70) <= packet_in;
						counter <= "0000010001011011";
						WHEN "0000010001011011" =>
						DD(11, 71) <= packet_in;
						counter <= "0000010001011100";
						WHEN "0000010001011100" =>
						DD(11, 72) <= packet_in;
						counter <= "0000010001011101";
						WHEN "0000010001011101" =>
						DD(11, 73) <= packet_in;
						counter <= "0000010001011110";
						WHEN "0000010001011110" =>
						DD(11, 74) <= packet_in;
						counter <= "0000010001011111";
						WHEN "0000010001011111" =>
						DD(11, 75) <= packet_in;
						counter <= "0000010001100000";
						WHEN "0000010001100000" =>
						DD(11, 76) <= packet_in;
						counter <= "0000010001100001";
						WHEN "0000010001100001" =>
						DD(11, 77) <= packet_in;
						counter <= "0000010001100010";
						WHEN "0000010001100010" =>
						DD(11, 78) <= packet_in;
						counter <= "0000010001100011";
						WHEN "0000010001100011" =>
						DD(11, 79) <= packet_in;
						counter <= "0000010001100100";
						WHEN "0000010001100100" =>
						DD(11, 80) <= packet_in;
						counter <= "0000010001100101";
						WHEN "0000010001100101" =>
						DD(11, 81) <= packet_in;
						counter <= "0000010001100110";
						WHEN "0000010001100110" =>
						DD(11, 82) <= packet_in;
						counter <= "0000010001100111";
						WHEN "0000010001100111" =>
						DD(11, 83) <= packet_in;
						counter <= "0000010001101000";
						WHEN "0000010001101000" =>
						DD(11, 84) <= packet_in;
						counter <= "0000010001101001";
						WHEN "0000010001101001" =>
						DD(11, 85) <= packet_in;
						counter <= "0000010001101010";
						WHEN "0000010001101010" =>
						DD(11, 86) <= packet_in;
						counter <= "0000010001101011";
						WHEN "0000010001101011" =>
						DD(11, 87) <= packet_in;
						counter <= "0000010001101100";
						WHEN "0000010001101100" =>
						DD(11, 88) <= packet_in;
						counter <= "0000010001101101";
						WHEN "0000010001101101" =>
						DD(11, 89) <= packet_in;
						counter <= "0000010001101110";
						WHEN "0000010001101110" =>
						DD(11, 90) <= packet_in;
						counter <= "0000010001101111";
						WHEN "0000010001101111" =>
						DD(11, 91) <= packet_in;
						counter <= "0000010001110000";
						WHEN "0000010001110000" =>
						DD(12, 0) <= packet_in;
						counter <= "0000010001110001";
						WHEN "0000010001110001" =>
						DD(12, 1) <= packet_in;
						counter <= "0000010001110010";
						WHEN "0000010001110010" =>
						DD(12, 2) <= packet_in;
						counter <= "0000010001110011";
						WHEN "0000010001110011" =>
						DD(12, 3) <= packet_in;
						counter <= "0000010001110100";
						WHEN "0000010001110100" =>
						DD(12, 4) <= packet_in;
						counter <= "0000010001110101";
						WHEN "0000010001110101" =>
						DD(12, 5) <= packet_in;
						counter <= "0000010001110110";
						WHEN "0000010001110110" =>
						DD(12, 6) <= packet_in;
						counter <= "0000010001110111";
						WHEN "0000010001110111" =>
						DD(12, 7) <= packet_in;
						counter <= "0000010001111000";
						WHEN "0000010001111000" =>
						DD(12, 8) <= packet_in;
						counter <= "0000010001111001";
						WHEN "0000010001111001" =>
						DD(12, 9) <= packet_in;
						counter <= "0000010001111010";
						WHEN "0000010001111010" =>
						DD(12, 10) <= packet_in;
						counter <= "0000010001111011";
						WHEN "0000010001111011" =>
						DD(12, 11) <= packet_in;
						counter <= "0000010001111100";
						WHEN "0000010001111100" =>
						DD(12, 12) <= packet_in;
						counter <= "0000010001111101";
						WHEN "0000010001111101" =>
						DD(12, 13) <= packet_in;
						counter <= "0000010001111110";
						WHEN "0000010001111110" =>
						DD(12, 14) <= packet_in;
						counter <= "0000010001111111";
						WHEN "0000010001111111" =>
						DD(12, 15) <= packet_in;
						counter <= "0000010010000000";
						WHEN "0000010010000000" =>
						DD(12, 16) <= packet_in;
						counter <= "0000010010000001";
						WHEN "0000010010000001" =>
						DD(12, 17) <= packet_in;
						counter <= "0000010010000010";
						WHEN "0000010010000010" =>
						DD(12, 18) <= packet_in;
						counter <= "0000010010000011";
						WHEN "0000010010000011" =>
						DD(12, 19) <= packet_in;
						counter <= "0000010010000100";
						WHEN "0000010010000100" =>
						DD(12, 20) <= packet_in;
						counter <= "0000010010000101";
						WHEN "0000010010000101" =>
						DD(12, 21) <= packet_in;
						counter <= "0000010010000110";
						WHEN "0000010010000110" =>
						DD(12, 22) <= packet_in;
						counter <= "0000010010000111";
						WHEN "0000010010000111" =>
						DD(12, 23) <= packet_in;
						counter <= "0000010010001000";
						WHEN "0000010010001000" =>
						DD(12, 24) <= packet_in;
						counter <= "0000010010001001";
						WHEN "0000010010001001" =>
						DD(12, 25) <= packet_in;
						counter <= "0000010010001010";
						WHEN "0000010010001010" =>
						DD(12, 26) <= packet_in;
						counter <= "0000010010001011";
						WHEN "0000010010001011" =>
						DD(12, 27) <= packet_in;
						counter <= "0000010010001100";
						WHEN "0000010010001100" =>
						DD(12, 28) <= packet_in;
						counter <= "0000010010001101";
						WHEN "0000010010001101" =>
						DD(12, 29) <= packet_in;
						counter <= "0000010010001110";
						WHEN "0000010010001110" =>
						DD(12, 30) <= packet_in;
						counter <= "0000010010001111";
						WHEN "0000010010001111" =>
						DD(12, 31) <= packet_in;
						counter <= "0000010010010000";
						WHEN "0000010010010000" =>
						DD(12, 32) <= packet_in;
						counter <= "0000010010010001";
						WHEN "0000010010010001" =>
						DD(12, 33) <= packet_in;
						counter <= "0000010010010010";
						WHEN "0000010010010010" =>
						DD(12, 34) <= packet_in;
						counter <= "0000010010010011";
						WHEN "0000010010010011" =>
						DD(12, 35) <= packet_in;
						counter <= "0000010010010100";
						WHEN "0000010010010100" =>
						DD(12, 36) <= packet_in;
						counter <= "0000010010010101";
						WHEN "0000010010010101" =>
						DD(12, 37) <= packet_in;
						counter <= "0000010010010110";
						WHEN "0000010010010110" =>
						DD(12, 38) <= packet_in;
						counter <= "0000010010010111";
						WHEN "0000010010010111" =>
						DD(12, 39) <= packet_in;
						counter <= "0000010010011000";
						WHEN "0000010010011000" =>
						DD(12, 40) <= packet_in;
						counter <= "0000010010011001";
						WHEN "0000010010011001" =>
						DD(12, 41) <= packet_in;
						counter <= "0000010010011010";
						WHEN "0000010010011010" =>
						DD(12, 42) <= packet_in;
						counter <= "0000010010011011";
						WHEN "0000010010011011" =>
						DD(12, 43) <= packet_in;
						counter <= "0000010010011100";
						WHEN "0000010010011100" =>
						DD(12, 44) <= packet_in;
						counter <= "0000010010011101";
						WHEN "0000010010011101" =>
						DD(12, 45) <= packet_in;
						counter <= "0000010010011110";
						WHEN "0000010010011110" =>
						DD(12, 46) <= packet_in;
						counter <= "0000010010011111";
						WHEN "0000010010011111" =>
						DD(12, 47) <= packet_in;
						counter <= "0000010010100000";
						WHEN "0000010010100000" =>
						DD(12, 48) <= packet_in;
						counter <= "0000010010100001";
						WHEN "0000010010100001" =>
						DD(12, 49) <= packet_in;
						counter <= "0000010010100010";
						WHEN "0000010010100010" =>
						DD(12, 50) <= packet_in;
						counter <= "0000010010100011";
						WHEN "0000010010100011" =>
						DD(12, 51) <= packet_in;
						counter <= "0000010010100100";
						WHEN "0000010010100100" =>
						DD(12, 52) <= packet_in;
						counter <= "0000010010100101";
						WHEN "0000010010100101" =>
						DD(12, 53) <= packet_in;
						counter <= "0000010010100110";
						WHEN "0000010010100110" =>
						DD(12, 54) <= packet_in;
						counter <= "0000010010100111";
						WHEN "0000010010100111" =>
						DD(12, 55) <= packet_in;
						counter <= "0000010010101000";
						WHEN "0000010010101000" =>
						DD(12, 56) <= packet_in;
						counter <= "0000010010101001";
						WHEN "0000010010101001" =>
						DD(12, 57) <= packet_in;
						counter <= "0000010010101010";
						WHEN "0000010010101010" =>
						DD(12, 58) <= packet_in;
						counter <= "0000010010101011";
						WHEN "0000010010101011" =>
						DD(12, 59) <= packet_in;
						counter <= "0000010010101100";
						WHEN "0000010010101100" =>
						DD(12, 60) <= packet_in;
						counter <= "0000010010101101";
						WHEN "0000010010101101" =>
						DD(12, 61) <= packet_in;
						counter <= "0000010010101110";
						WHEN "0000010010101110" =>
						DD(12, 62) <= packet_in;
						counter <= "0000010010101111";
						WHEN "0000010010101111" =>
						DD(12, 63) <= packet_in;
						counter <= "0000010010110000";
						WHEN "0000010010110000" =>
						DD(12, 64) <= packet_in;
						counter <= "0000010010110001";
						WHEN "0000010010110001" =>
						DD(12, 65) <= packet_in;
						counter <= "0000010010110010";
						WHEN "0000010010110010" =>
						DD(12, 66) <= packet_in;
						counter <= "0000010010110011";
						WHEN "0000010010110011" =>
						DD(12, 67) <= packet_in;
						counter <= "0000010010110100";
						WHEN "0000010010110100" =>
						DD(12, 68) <= packet_in;
						counter <= "0000010010110101";
						WHEN "0000010010110101" =>
						DD(12, 69) <= packet_in;
						counter <= "0000010010110110";
						WHEN "0000010010110110" =>
						DD(12, 70) <= packet_in;
						counter <= "0000010010110111";
						WHEN "0000010010110111" =>
						DD(12, 71) <= packet_in;
						counter <= "0000010010111000";
						WHEN "0000010010111000" =>
						DD(12, 72) <= packet_in;
						counter <= "0000010010111001";
						WHEN "0000010010111001" =>
						DD(12, 73) <= packet_in;
						counter <= "0000010010111010";
						WHEN "0000010010111010" =>
						DD(12, 74) <= packet_in;
						counter <= "0000010010111011";
						WHEN "0000010010111011" =>
						DD(12, 75) <= packet_in;
						counter <= "0000010010111100";
						WHEN "0000010010111100" =>
						DD(12, 76) <= packet_in;
						counter <= "0000010010111101";
						WHEN "0000010010111101" =>
						DD(12, 77) <= packet_in;
						counter <= "0000010010111110";
						WHEN "0000010010111110" =>
						DD(12, 78) <= packet_in;
						counter <= "0000010010111111";
						WHEN "0000010010111111" =>
						DD(12, 79) <= packet_in;
						counter <= "0000010011000000";
						WHEN "0000010011000000" =>
						DD(12, 80) <= packet_in;
						counter <= "0000010011000001";
						WHEN "0000010011000001" =>
						DD(12, 81) <= packet_in;
						counter <= "0000010011000010";
						WHEN "0000010011000010" =>
						DD(12, 82) <= packet_in;
						counter <= "0000010011000011";
						WHEN "0000010011000011" =>
						DD(12, 83) <= packet_in;
						counter <= "0000010011000100";
						WHEN "0000010011000100" =>
						DD(12, 84) <= packet_in;
						counter <= "0000010011000101";
						WHEN "0000010011000101" =>
						DD(12, 85) <= packet_in;
						counter <= "0000010011000110";
						WHEN "0000010011000110" =>
						DD(12, 86) <= packet_in;
						counter <= "0000010011000111";
						WHEN "0000010011000111" =>
						DD(12, 87) <= packet_in;
						counter <= "0000010011001000";
						WHEN "0000010011001000" =>
						DD(12, 88) <= packet_in;
						counter <= "0000010011001001";
						WHEN "0000010011001001" =>
						DD(12, 89) <= packet_in;
						counter <= "0000010011001010";
						WHEN "0000010011001010" =>
						DD(12, 90) <= packet_in;
						counter <= "0000010011001011";
						WHEN "0000010011001011" =>
						DD(12, 91) <= packet_in;
						counter <= "0000010011001100";
						WHEN "0000010011001100" =>
						DD(13, 0) <= packet_in;
						counter <= "0000010011001101";
						WHEN "0000010011001101" =>
						DD(13, 1) <= packet_in;
						counter <= "0000010011001110";
						WHEN "0000010011001110" =>
						DD(13, 2) <= packet_in;
						counter <= "0000010011001111";
						WHEN "0000010011001111" =>
						DD(13, 3) <= packet_in;
						counter <= "0000010011010000";
						WHEN "0000010011010000" =>
						DD(13, 4) <= packet_in;
						counter <= "0000010011010001";
						WHEN "0000010011010001" =>
						DD(13, 5) <= packet_in;
						counter <= "0000010011010010";
						WHEN "0000010011010010" =>
						DD(13, 6) <= packet_in;
						counter <= "0000010011010011";
						WHEN "0000010011010011" =>
						DD(13, 7) <= packet_in;
						counter <= "0000010011010100";
						WHEN "0000010011010100" =>
						DD(13, 8) <= packet_in;
						counter <= "0000010011010101";
						WHEN "0000010011010101" =>
						DD(13, 9) <= packet_in;
						counter <= "0000010011010110";
						WHEN "0000010011010110" =>
						DD(13, 10) <= packet_in;
						counter <= "0000010011010111";
						WHEN "0000010011010111" =>
						DD(13, 11) <= packet_in;
						counter <= "0000010011011000";
						WHEN "0000010011011000" =>
						DD(13, 12) <= packet_in;
						counter <= "0000010011011001";
						WHEN "0000010011011001" =>
						DD(13, 13) <= packet_in;
						counter <= "0000010011011010";
						WHEN "0000010011011010" =>
						DD(13, 14) <= packet_in;
						counter <= "0000010011011011";
						WHEN "0000010011011011" =>
						DD(13, 15) <= packet_in;
						counter <= "0000010011011100";
						WHEN "0000010011011100" =>
						DD(13, 16) <= packet_in;
						counter <= "0000010011011101";
						WHEN "0000010011011101" =>
						DD(13, 17) <= packet_in;
						counter <= "0000010011011110";
						WHEN "0000010011011110" =>
						DD(13, 18) <= packet_in;
						counter <= "0000010011011111";
						WHEN "0000010011011111" =>
						DD(13, 19) <= packet_in;
						counter <= "0000010011100000";
						WHEN "0000010011100000" =>
						DD(13, 20) <= packet_in;
						counter <= "0000010011100001";
						WHEN "0000010011100001" =>
						DD(13, 21) <= packet_in;
						counter <= "0000010011100010";
						WHEN "0000010011100010" =>
						DD(13, 22) <= packet_in;
						counter <= "0000010011100011";
						WHEN "0000010011100011" =>
						DD(13, 23) <= packet_in;
						counter <= "0000010011100100";
						WHEN "0000010011100100" =>
						DD(13, 24) <= packet_in;
						counter <= "0000010011100101";
						WHEN "0000010011100101" =>
						DD(13, 25) <= packet_in;
						counter <= "0000010011100110";
						WHEN "0000010011100110" =>
						DD(13, 26) <= packet_in;
						counter <= "0000010011100111";
						WHEN "0000010011100111" =>
						DD(13, 27) <= packet_in;
						counter <= "0000010011101000";
						WHEN "0000010011101000" =>
						DD(13, 28) <= packet_in;
						counter <= "0000010011101001";
						WHEN "0000010011101001" =>
						DD(13, 29) <= packet_in;
						counter <= "0000010011101010";
						WHEN "0000010011101010" =>
						DD(13, 30) <= packet_in;
						counter <= "0000010011101011";
						WHEN "0000010011101011" =>
						DD(13, 31) <= packet_in;
						counter <= "0000010011101100";
						WHEN "0000010011101100" =>
						DD(13, 32) <= packet_in;
						counter <= "0000010011101101";
						WHEN "0000010011101101" =>
						DD(13, 33) <= packet_in;
						counter <= "0000010011101110";
						WHEN "0000010011101110" =>
						DD(13, 34) <= packet_in;
						counter <= "0000010011101111";
						WHEN "0000010011101111" =>
						DD(13, 35) <= packet_in;
						counter <= "0000010011110000";
						WHEN "0000010011110000" =>
						DD(13, 36) <= packet_in;
						counter <= "0000010011110001";
						WHEN "0000010011110001" =>
						DD(13, 37) <= packet_in;
						counter <= "0000010011110010";
						WHEN "0000010011110010" =>
						DD(13, 38) <= packet_in;
						counter <= "0000010011110011";
						WHEN "0000010011110011" =>
						DD(13, 39) <= packet_in;
						counter <= "0000010011110100";
						WHEN "0000010011110100" =>
						DD(13, 40) <= packet_in;
						counter <= "0000010011110101";
						WHEN "0000010011110101" =>
						DD(13, 41) <= packet_in;
						counter <= "0000010011110110";
						WHEN "0000010011110110" =>
						DD(13, 42) <= packet_in;
						counter <= "0000010011110111";
						WHEN "0000010011110111" =>
						DD(13, 43) <= packet_in;
						counter <= "0000010011111000";
						WHEN "0000010011111000" =>
						DD(13, 44) <= packet_in;
						counter <= "0000010011111001";
						WHEN "0000010011111001" =>
						DD(13, 45) <= packet_in;
						counter <= "0000010011111010";
						WHEN "0000010011111010" =>
						DD(13, 46) <= packet_in;
						counter <= "0000010011111011";
						WHEN "0000010011111011" =>
						DD(13, 47) <= packet_in;
						counter <= "0000010011111100";
						WHEN "0000010011111100" =>
						DD(13, 48) <= packet_in;
						counter <= "0000010011111101";
						WHEN "0000010011111101" =>
						DD(13, 49) <= packet_in;
						counter <= "0000010011111110";
						WHEN "0000010011111110" =>
						DD(13, 50) <= packet_in;
						counter <= "0000010011111111";
						WHEN "0000010011111111" =>
						DD(13, 51) <= packet_in;
						counter <= "0000010100000000";
						WHEN "0000010100000000" =>
						DD(13, 52) <= packet_in;
						counter <= "0000010100000001";
						WHEN "0000010100000001" =>
						DD(13, 53) <= packet_in;
						counter <= "0000010100000010";
						WHEN "0000010100000010" =>
						DD(13, 54) <= packet_in;
						counter <= "0000010100000011";
						WHEN "0000010100000011" =>
						DD(13, 55) <= packet_in;
						counter <= "0000010100000100";
						WHEN "0000010100000100" =>
						DD(13, 56) <= packet_in;
						counter <= "0000010100000101";
						WHEN "0000010100000101" =>
						DD(13, 57) <= packet_in;
						counter <= "0000010100000110";
						WHEN "0000010100000110" =>
						DD(13, 58) <= packet_in;
						counter <= "0000010100000111";
						WHEN "0000010100000111" =>
						DD(13, 59) <= packet_in;
						counter <= "0000010100001000";
						WHEN "0000010100001000" =>
						DD(13, 60) <= packet_in;
						counter <= "0000010100001001";
						WHEN "0000010100001001" =>
						DD(13, 61) <= packet_in;
						counter <= "0000010100001010";
						WHEN "0000010100001010" =>
						DD(13, 62) <= packet_in;
						counter <= "0000010100001011";
						WHEN "0000010100001011" =>
						DD(13, 63) <= packet_in;
						counter <= "0000010100001100";
						WHEN "0000010100001100" =>
						DD(13, 64) <= packet_in;
						counter <= "0000010100001101";
						WHEN "0000010100001101" =>
						DD(13, 65) <= packet_in;
						counter <= "0000010100001110";
						WHEN "0000010100001110" =>
						DD(13, 66) <= packet_in;
						counter <= "0000010100001111";
						WHEN "0000010100001111" =>
						DD(13, 67) <= packet_in;
						counter <= "0000010100010000";
						WHEN "0000010100010000" =>
						DD(13, 68) <= packet_in;
						counter <= "0000010100010001";
						WHEN "0000010100010001" =>
						DD(13, 69) <= packet_in;
						counter <= "0000010100010010";
						WHEN "0000010100010010" =>
						DD(13, 70) <= packet_in;
						counter <= "0000010100010011";
						WHEN "0000010100010011" =>
						DD(13, 71) <= packet_in;
						counter <= "0000010100010100";
						WHEN "0000010100010100" =>
						DD(13, 72) <= packet_in;
						counter <= "0000010100010101";
						WHEN "0000010100010101" =>
						DD(13, 73) <= packet_in;
						counter <= "0000010100010110";
						WHEN "0000010100010110" =>
						DD(13, 74) <= packet_in;
						counter <= "0000010100010111";
						WHEN "0000010100010111" =>
						DD(13, 75) <= packet_in;
						counter <= "0000010100011000";
						WHEN "0000010100011000" =>
						DD(13, 76) <= packet_in;
						counter <= "0000010100011001";
						WHEN "0000010100011001" =>
						DD(13, 77) <= packet_in;
						counter <= "0000010100011010";
						WHEN "0000010100011010" =>
						DD(13, 78) <= packet_in;
						counter <= "0000010100011011";
						WHEN "0000010100011011" =>
						DD(13, 79) <= packet_in;
						counter <= "0000010100011100";
						WHEN "0000010100011100" =>
						DD(13, 80) <= packet_in;
						counter <= "0000010100011101";
						WHEN "0000010100011101" =>
						DD(13, 81) <= packet_in;
						counter <= "0000010100011110";
						WHEN "0000010100011110" =>
						DD(13, 82) <= packet_in;
						counter <= "0000010100011111";
						WHEN "0000010100011111" =>
						DD(13, 83) <= packet_in;
						counter <= "0000010100100000";
						WHEN "0000010100100000" =>
						DD(13, 84) <= packet_in;
						counter <= "0000010100100001";
						WHEN "0000010100100001" =>
						DD(13, 85) <= packet_in;
						counter <= "0000010100100010";
						WHEN "0000010100100010" =>
						DD(13, 86) <= packet_in;
						counter <= "0000010100100011";
						WHEN "0000010100100011" =>
						DD(13, 87) <= packet_in;
						counter <= "0000010100100100";
						WHEN "0000010100100100" =>
						DD(13, 88) <= packet_in;
						counter <= "0000010100100101";
						WHEN "0000010100100101" =>
						DD(13, 89) <= packet_in;
						counter <= "0000010100100110";
						WHEN "0000010100100110" =>
						DD(13, 90) <= packet_in;
						counter <= "0000010100100111";
						WHEN "0000010100100111" =>
						DD(13, 91) <= packet_in;
						counter <= "0000010100101000";
						WHEN "0000010100101000" =>
						DD(14, 0) <= packet_in;
						counter <= "0000010100101001";
						WHEN "0000010100101001" =>
						DD(14, 1) <= packet_in;
						counter <= "0000010100101010";
						WHEN "0000010100101010" =>
						DD(14, 2) <= packet_in;
						counter <= "0000010100101011";
						WHEN "0000010100101011" =>
						DD(14, 3) <= packet_in;
						counter <= "0000010100101100";
						WHEN "0000010100101100" =>
						DD(14, 4) <= packet_in;
						counter <= "0000010100101101";
						WHEN "0000010100101101" =>
						DD(14, 5) <= packet_in;
						counter <= "0000010100101110";
						WHEN "0000010100101110" =>
						DD(14, 6) <= packet_in;
						counter <= "0000010100101111";
						WHEN "0000010100101111" =>
						DD(14, 7) <= packet_in;
						counter <= "0000010100110000";
						WHEN "0000010100110000" =>
						DD(14, 8) <= packet_in;
						counter <= "0000010100110001";
						WHEN "0000010100110001" =>
						DD(14, 9) <= packet_in;
						counter <= "0000010100110010";
						WHEN "0000010100110010" =>
						DD(14, 10) <= packet_in;
						counter <= "0000010100110011";
						WHEN "0000010100110011" =>
						DD(14, 11) <= packet_in;
						counter <= "0000010100110100";
						WHEN "0000010100110100" =>
						DD(14, 12) <= packet_in;
						counter <= "0000010100110101";
						WHEN "0000010100110101" =>
						DD(14, 13) <= packet_in;
						counter <= "0000010100110110";
						WHEN "0000010100110110" =>
						DD(14, 14) <= packet_in;
						counter <= "0000010100110111";
						WHEN "0000010100110111" =>
						DD(14, 15) <= packet_in;
						counter <= "0000010100111000";
						WHEN "0000010100111000" =>
						DD(14, 16) <= packet_in;
						counter <= "0000010100111001";
						WHEN "0000010100111001" =>
						DD(14, 17) <= packet_in;
						counter <= "0000010100111010";
						WHEN "0000010100111010" =>
						DD(14, 18) <= packet_in;
						counter <= "0000010100111011";
						WHEN "0000010100111011" =>
						DD(14, 19) <= packet_in;
						counter <= "0000010100111100";
						WHEN "0000010100111100" =>
						DD(14, 20) <= packet_in;
						counter <= "0000010100111101";
						WHEN "0000010100111101" =>
						DD(14, 21) <= packet_in;
						counter <= "0000010100111110";
						WHEN "0000010100111110" =>
						DD(14, 22) <= packet_in;
						counter <= "0000010100111111";
						WHEN "0000010100111111" =>
						DD(14, 23) <= packet_in;
						counter <= "0000010101000000";
						WHEN "0000010101000000" =>
						DD(14, 24) <= packet_in;
						counter <= "0000010101000001";
						WHEN "0000010101000001" =>
						DD(14, 25) <= packet_in;
						counter <= "0000010101000010";
						WHEN "0000010101000010" =>
						DD(14, 26) <= packet_in;
						counter <= "0000010101000011";
						WHEN "0000010101000011" =>
						DD(14, 27) <= packet_in;
						counter <= "0000010101000100";
						WHEN "0000010101000100" =>
						DD(14, 28) <= packet_in;
						counter <= "0000010101000101";
						WHEN "0000010101000101" =>
						DD(14, 29) <= packet_in;
						counter <= "0000010101000110";
						WHEN "0000010101000110" =>
						DD(14, 30) <= packet_in;
						counter <= "0000010101000111";
						WHEN "0000010101000111" =>
						DD(14, 31) <= packet_in;
						counter <= "0000010101001000";
						WHEN "0000010101001000" =>
						DD(14, 32) <= packet_in;
						counter <= "0000010101001001";
						WHEN "0000010101001001" =>
						DD(14, 33) <= packet_in;
						counter <= "0000010101001010";
						WHEN "0000010101001010" =>
						DD(14, 34) <= packet_in;
						counter <= "0000010101001011";
						WHEN "0000010101001011" =>
						DD(14, 35) <= packet_in;
						counter <= "0000010101001100";
						WHEN "0000010101001100" =>
						DD(14, 36) <= packet_in;
						counter <= "0000010101001101";
						WHEN "0000010101001101" =>
						DD(14, 37) <= packet_in;
						counter <= "0000010101001110";
						WHEN "0000010101001110" =>
						DD(14, 38) <= packet_in;
						counter <= "0000010101001111";
						WHEN "0000010101001111" =>
						DD(14, 39) <= packet_in;
						counter <= "0000010101010000";
						WHEN "0000010101010000" =>
						DD(14, 40) <= packet_in;
						counter <= "0000010101010001";
						WHEN "0000010101010001" =>
						DD(14, 41) <= packet_in;
						counter <= "0000010101010010";
						WHEN "0000010101010010" =>
						DD(14, 42) <= packet_in;
						counter <= "0000010101010011";
						WHEN "0000010101010011" =>
						DD(14, 43) <= packet_in;
						counter <= "0000010101010100";
						WHEN "0000010101010100" =>
						DD(14, 44) <= packet_in;
						counter <= "0000010101010101";
						WHEN "0000010101010101" =>
						DD(14, 45) <= packet_in;
						counter <= "0000010101010110";
						WHEN "0000010101010110" =>
						DD(14, 46) <= packet_in;
						counter <= "0000010101010111";
						WHEN "0000010101010111" =>
						DD(14, 47) <= packet_in;
						counter <= "0000010101011000";
						WHEN "0000010101011000" =>
						DD(14, 48) <= packet_in;
						counter <= "0000010101011001";
						WHEN "0000010101011001" =>
						DD(14, 49) <= packet_in;
						counter <= "0000010101011010";
						WHEN "0000010101011010" =>
						DD(14, 50) <= packet_in;
						counter <= "0000010101011011";
						WHEN "0000010101011011" =>
						DD(14, 51) <= packet_in;
						counter <= "0000010101011100";
						WHEN "0000010101011100" =>
						DD(14, 52) <= packet_in;
						counter <= "0000010101011101";
						WHEN "0000010101011101" =>
						DD(14, 53) <= packet_in;
						counter <= "0000010101011110";
						WHEN "0000010101011110" =>
						DD(14, 54) <= packet_in;
						counter <= "0000010101011111";
						WHEN "0000010101011111" =>
						DD(14, 55) <= packet_in;
						counter <= "0000010101100000";
						WHEN "0000010101100000" =>
						DD(14, 56) <= packet_in;
						counter <= "0000010101100001";
						WHEN "0000010101100001" =>
						DD(14, 57) <= packet_in;
						counter <= "0000010101100010";
						WHEN "0000010101100010" =>
						DD(14, 58) <= packet_in;
						counter <= "0000010101100011";
						WHEN "0000010101100011" =>
						DD(14, 59) <= packet_in;
						counter <= "0000010101100100";
						WHEN "0000010101100100" =>
						DD(14, 60) <= packet_in;
						counter <= "0000010101100101";
						WHEN "0000010101100101" =>
						DD(14, 61) <= packet_in;
						counter <= "0000010101100110";
						WHEN "0000010101100110" =>
						DD(14, 62) <= packet_in;
						counter <= "0000010101100111";
						WHEN "0000010101100111" =>
						DD(14, 63) <= packet_in;
						counter <= "0000010101101000";
						WHEN "0000010101101000" =>
						DD(14, 64) <= packet_in;
						counter <= "0000010101101001";
						WHEN "0000010101101001" =>
						DD(14, 65) <= packet_in;
						counter <= "0000010101101010";
						WHEN "0000010101101010" =>
						DD(14, 66) <= packet_in;
						counter <= "0000010101101011";
						WHEN "0000010101101011" =>
						DD(14, 67) <= packet_in;
						counter <= "0000010101101100";
						WHEN "0000010101101100" =>
						DD(14, 68) <= packet_in;
						counter <= "0000010101101101";
						WHEN "0000010101101101" =>
						DD(14, 69) <= packet_in;
						counter <= "0000010101101110";
						WHEN "0000010101101110" =>
						DD(14, 70) <= packet_in;
						counter <= "0000010101101111";
						WHEN "0000010101101111" =>
						DD(14, 71) <= packet_in;
						counter <= "0000010101110000";
						WHEN "0000010101110000" =>
						DD(14, 72) <= packet_in;
						counter <= "0000010101110001";
						WHEN "0000010101110001" =>
						DD(14, 73) <= packet_in;
						counter <= "0000010101110010";
						WHEN "0000010101110010" =>
						DD(14, 74) <= packet_in;
						counter <= "0000010101110011";
						WHEN "0000010101110011" =>
						DD(14, 75) <= packet_in;
						counter <= "0000010101110100";
						WHEN "0000010101110100" =>
						DD(14, 76) <= packet_in;
						counter <= "0000010101110101";
						WHEN "0000010101110101" =>
						DD(14, 77) <= packet_in;
						counter <= "0000010101110110";
						WHEN "0000010101110110" =>
						DD(14, 78) <= packet_in;
						counter <= "0000010101110111";
						WHEN "0000010101110111" =>
						DD(14, 79) <= packet_in;
						counter <= "0000010101111000";
						WHEN "0000010101111000" =>
						DD(14, 80) <= packet_in;
						counter <= "0000010101111001";
						WHEN "0000010101111001" =>
						DD(14, 81) <= packet_in;
						counter <= "0000010101111010";
						WHEN "0000010101111010" =>
						DD(14, 82) <= packet_in;
						counter <= "0000010101111011";
						WHEN "0000010101111011" =>
						DD(14, 83) <= packet_in;
						counter <= "0000010101111100";
						WHEN "0000010101111100" =>
						DD(14, 84) <= packet_in;
						counter <= "0000010101111101";
						WHEN "0000010101111101" =>
						DD(14, 85) <= packet_in;
						counter <= "0000010101111110";
						WHEN "0000010101111110" =>
						DD(14, 86) <= packet_in;
						counter <= "0000010101111111";
						WHEN "0000010101111111" =>
						DD(14, 87) <= packet_in;
						counter <= "0000010110000000";
						WHEN "0000010110000000" =>
						DD(14, 88) <= packet_in;
						counter <= "0000010110000001";
						WHEN "0000010110000001" =>
						DD(14, 89) <= packet_in;
						counter <= "0000010110000010";
						WHEN "0000010110000010" =>
						DD(14, 90) <= packet_in;
						counter <= "0000010110000011";
						WHEN "0000010110000011" =>
						DD(14, 91) <= packet_in;
						counter <= "0000010110000100";
						WHEN "0000010110000100" =>
						DD(15, 0) <= packet_in;
						counter <= "0000010110000101";
						WHEN "0000010110000101" =>
						DD(15, 1) <= packet_in;
						counter <= "0000010110000110";
						WHEN "0000010110000110" =>
						DD(15, 2) <= packet_in;
						counter <= "0000010110000111";
						WHEN "0000010110000111" =>
						DD(15, 3) <= packet_in;
						counter <= "0000010110001000";
						WHEN "0000010110001000" =>
						DD(15, 4) <= packet_in;
						counter <= "0000010110001001";
						WHEN "0000010110001001" =>
						DD(15, 5) <= packet_in;
						counter <= "0000010110001010";
						WHEN "0000010110001010" =>
						DD(15, 6) <= packet_in;
						counter <= "0000010110001011";
						WHEN "0000010110001011" =>
						DD(15, 7) <= packet_in;
						counter <= "0000010110001100";
						WHEN "0000010110001100" =>
						DD(15, 8) <= packet_in;
						counter <= "0000010110001101";
						WHEN "0000010110001101" =>
						DD(15, 9) <= packet_in;
						counter <= "0000010110001110";
						WHEN "0000010110001110" =>
						DD(15, 10) <= packet_in;
						counter <= "0000010110001111";
						WHEN "0000010110001111" =>
						DD(15, 11) <= packet_in;
						counter <= "0000010110010000";
						WHEN "0000010110010000" =>
						DD(15, 12) <= packet_in;
						counter <= "0000010110010001";
						WHEN "0000010110010001" =>
						DD(15, 13) <= packet_in;
						counter <= "0000010110010010";
						WHEN "0000010110010010" =>
						DD(15, 14) <= packet_in;
						counter <= "0000010110010011";
						WHEN "0000010110010011" =>
						DD(15, 15) <= packet_in;
						counter <= "0000010110010100";
						WHEN "0000010110010100" =>
						DD(15, 16) <= packet_in;
						counter <= "0000010110010101";
						WHEN "0000010110010101" =>
						DD(15, 17) <= packet_in;
						counter <= "0000010110010110";
						WHEN "0000010110010110" =>
						DD(15, 18) <= packet_in;
						counter <= "0000010110010111";
						WHEN "0000010110010111" =>
						DD(15, 19) <= packet_in;
						counter <= "0000010110011000";
						WHEN "0000010110011000" =>
						DD(15, 20) <= packet_in;
						counter <= "0000010110011001";
						WHEN "0000010110011001" =>
						DD(15, 21) <= packet_in;
						counter <= "0000010110011010";
						WHEN "0000010110011010" =>
						DD(15, 22) <= packet_in;
						counter <= "0000010110011011";
						WHEN "0000010110011011" =>
						DD(15, 23) <= packet_in;
						counter <= "0000010110011100";
						WHEN "0000010110011100" =>
						DD(15, 24) <= packet_in;
						counter <= "0000010110011101";
						WHEN "0000010110011101" =>
						DD(15, 25) <= packet_in;
						counter <= "0000010110011110";
						WHEN "0000010110011110" =>
						DD(15, 26) <= packet_in;
						counter <= "0000010110011111";
						WHEN "0000010110011111" =>
						DD(15, 27) <= packet_in;
						counter <= "0000010110100000";
						WHEN "0000010110100000" =>
						DD(15, 28) <= packet_in;
						counter <= "0000010110100001";
						WHEN "0000010110100001" =>
						DD(15, 29) <= packet_in;
						counter <= "0000010110100010";
						WHEN "0000010110100010" =>
						DD(15, 30) <= packet_in;
						counter <= "0000010110100011";
						WHEN "0000010110100011" =>
						DD(15, 31) <= packet_in;
						counter <= "0000010110100100";
						WHEN "0000010110100100" =>
						DD(15, 32) <= packet_in;
						counter <= "0000010110100101";
						WHEN "0000010110100101" =>
						DD(15, 33) <= packet_in;
						counter <= "0000010110100110";
						WHEN "0000010110100110" =>
						DD(15, 34) <= packet_in;
						counter <= "0000010110100111";
						WHEN "0000010110100111" =>
						DD(15, 35) <= packet_in;
						counter <= "0000010110101000";
						WHEN "0000010110101000" =>
						DD(15, 36) <= packet_in;
						counter <= "0000010110101001";
						WHEN "0000010110101001" =>
						DD(15, 37) <= packet_in;
						counter <= "0000010110101010";
						WHEN "0000010110101010" =>
						DD(15, 38) <= packet_in;
						counter <= "0000010110101011";
						WHEN "0000010110101011" =>
						DD(15, 39) <= packet_in;
						counter <= "0000010110101100";
						WHEN "0000010110101100" =>
						DD(15, 40) <= packet_in;
						counter <= "0000010110101101";
						WHEN "0000010110101101" =>
						DD(15, 41) <= packet_in;
						counter <= "0000010110101110";
						WHEN "0000010110101110" =>
						DD(15, 42) <= packet_in;
						counter <= "0000010110101111";
						WHEN "0000010110101111" =>
						DD(15, 43) <= packet_in;
						counter <= "0000010110110000";
						WHEN "0000010110110000" =>
						DD(15, 44) <= packet_in;
						counter <= "0000010110110001";
						WHEN "0000010110110001" =>
						DD(15, 45) <= packet_in;
						counter <= "0000010110110010";
						WHEN "0000010110110010" =>
						DD(15, 46) <= packet_in;
						counter <= "0000010110110011";
						WHEN "0000010110110011" =>
						DD(15, 47) <= packet_in;
						counter <= "0000010110110100";
						WHEN "0000010110110100" =>
						DD(15, 48) <= packet_in;
						counter <= "0000010110110101";
						WHEN "0000010110110101" =>
						DD(15, 49) <= packet_in;
						counter <= "0000010110110110";
						WHEN "0000010110110110" =>
						DD(15, 50) <= packet_in;
						counter <= "0000010110110111";
						WHEN "0000010110110111" =>
						DD(15, 51) <= packet_in;
						counter <= "0000010110111000";
						WHEN "0000010110111000" =>
						DD(15, 52) <= packet_in;
						counter <= "0000010110111001";
						WHEN "0000010110111001" =>
						DD(15, 53) <= packet_in;
						counter <= "0000010110111010";
						WHEN "0000010110111010" =>
						DD(15, 54) <= packet_in;
						counter <= "0000010110111011";
						WHEN "0000010110111011" =>
						DD(15, 55) <= packet_in;
						counter <= "0000010110111100";
						WHEN "0000010110111100" =>
						DD(15, 56) <= packet_in;
						counter <= "0000010110111101";
						WHEN "0000010110111101" =>
						DD(15, 57) <= packet_in;
						counter <= "0000010110111110";
						WHEN "0000010110111110" =>
						DD(15, 58) <= packet_in;
						counter <= "0000010110111111";
						WHEN "0000010110111111" =>
						DD(15, 59) <= packet_in;
						counter <= "0000010111000000";
						WHEN "0000010111000000" =>
						DD(15, 60) <= packet_in;
						counter <= "0000010111000001";
						WHEN "0000010111000001" =>
						DD(15, 61) <= packet_in;
						counter <= "0000010111000010";
						WHEN "0000010111000010" =>
						DD(15, 62) <= packet_in;
						counter <= "0000010111000011";
						WHEN "0000010111000011" =>
						DD(15, 63) <= packet_in;
						counter <= "0000010111000100";
						WHEN "0000010111000100" =>
						DD(15, 64) <= packet_in;
						counter <= "0000010111000101";
						WHEN "0000010111000101" =>
						DD(15, 65) <= packet_in;
						counter <= "0000010111000110";
						WHEN "0000010111000110" =>
						DD(15, 66) <= packet_in;
						counter <= "0000010111000111";
						WHEN "0000010111000111" =>
						DD(15, 67) <= packet_in;
						counter <= "0000010111001000";
						WHEN "0000010111001000" =>
						DD(15, 68) <= packet_in;
						counter <= "0000010111001001";
						WHEN "0000010111001001" =>
						DD(15, 69) <= packet_in;
						counter <= "0000010111001010";
						WHEN "0000010111001010" =>
						DD(15, 70) <= packet_in;
						counter <= "0000010111001011";
						WHEN "0000010111001011" =>
						DD(15, 71) <= packet_in;
						counter <= "0000010111001100";
						WHEN "0000010111001100" =>
						DD(15, 72) <= packet_in;
						counter <= "0000010111001101";
						WHEN "0000010111001101" =>
						DD(15, 73) <= packet_in;
						counter <= "0000010111001110";
						WHEN "0000010111001110" =>
						DD(15, 74) <= packet_in;
						counter <= "0000010111001111";
						WHEN "0000010111001111" =>
						DD(15, 75) <= packet_in;
						counter <= "0000010111010000";
						WHEN "0000010111010000" =>
						DD(15, 76) <= packet_in;
						counter <= "0000010111010001";
						WHEN "0000010111010001" =>
						DD(15, 77) <= packet_in;
						counter <= "0000010111010010";
						WHEN "0000010111010010" =>
						DD(15, 78) <= packet_in;
						counter <= "0000010111010011";
						WHEN "0000010111010011" =>
						DD(15, 79) <= packet_in;
						counter <= "0000010111010100";
						WHEN "0000010111010100" =>
						DD(15, 80) <= packet_in;
						counter <= "0000010111010101";
						WHEN "0000010111010101" =>
						DD(15, 81) <= packet_in;
						counter <= "0000010111010110";
						WHEN "0000010111010110" =>
						DD(15, 82) <= packet_in;
						counter <= "0000010111010111";
						WHEN "0000010111010111" =>
						DD(15, 83) <= packet_in;
						counter <= "0000010111011000";
						WHEN "0000010111011000" =>
						DD(15, 84) <= packet_in;
						counter <= "0000010111011001";
						WHEN "0000010111011001" =>
						DD(15, 85) <= packet_in;
						counter <= "0000010111011010";
						WHEN "0000010111011010" =>
						DD(15, 86) <= packet_in;
						counter <= "0000010111011011";
						WHEN "0000010111011011" =>
						DD(15, 87) <= packet_in;
						counter <= "0000010111011100";
						WHEN "0000010111011100" =>
						DD(15, 88) <= packet_in;
						counter <= "0000010111011101";
						WHEN "0000010111011101" =>
						DD(15, 89) <= packet_in;
						counter <= "0000010111011110";
						WHEN "0000010111011110" =>
						DD(15, 90) <= packet_in;
						counter <= "0000010111011111";
						WHEN "0000010111011111" =>
						DD(15, 91) <= packet_in;
						counter <= "0000010111100000";
						WHEN "0000010111100000" =>
						DD(16, 0) <= packet_in;
						counter <= "0000010111100001";
						WHEN "0000010111100001" =>
						DD(16, 1) <= packet_in;
						counter <= "0000010111100010";
						WHEN "0000010111100010" =>
						DD(16, 2) <= packet_in;
						counter <= "0000010111100011";
						WHEN "0000010111100011" =>
						DD(16, 3) <= packet_in;
						counter <= "0000010111100100";
						WHEN "0000010111100100" =>
						DD(16, 4) <= packet_in;
						counter <= "0000010111100101";
						WHEN "0000010111100101" =>
						DD(16, 5) <= packet_in;
						counter <= "0000010111100110";
						WHEN "0000010111100110" =>
						DD(16, 6) <= packet_in;
						counter <= "0000010111100111";
						WHEN "0000010111100111" =>
						DD(16, 7) <= packet_in;
						counter <= "0000010111101000";
						WHEN "0000010111101000" =>
						DD(16, 8) <= packet_in;
						counter <= "0000010111101001";
						WHEN "0000010111101001" =>
						DD(16, 9) <= packet_in;
						counter <= "0000010111101010";
						WHEN "0000010111101010" =>
						DD(16, 10) <= packet_in;
						counter <= "0000010111101011";
						WHEN "0000010111101011" =>
						DD(16, 11) <= packet_in;
						counter <= "0000010111101100";
						WHEN "0000010111101100" =>
						DD(16, 12) <= packet_in;
						counter <= "0000010111101101";
						WHEN "0000010111101101" =>
						DD(16, 13) <= packet_in;
						counter <= "0000010111101110";
						WHEN "0000010111101110" =>
						DD(16, 14) <= packet_in;
						counter <= "0000010111101111";
						WHEN "0000010111101111" =>
						DD(16, 15) <= packet_in;
						counter <= "0000010111110000";
						WHEN "0000010111110000" =>
						DD(16, 16) <= packet_in;
						counter <= "0000010111110001";
						WHEN "0000010111110001" =>
						DD(16, 17) <= packet_in;
						counter <= "0000010111110010";
						WHEN "0000010111110010" =>
						DD(16, 18) <= packet_in;
						counter <= "0000010111110011";
						WHEN "0000010111110011" =>
						DD(16, 19) <= packet_in;
						counter <= "0000010111110100";
						WHEN "0000010111110100" =>
						DD(16, 20) <= packet_in;
						counter <= "0000010111110101";
						WHEN "0000010111110101" =>
						DD(16, 21) <= packet_in;
						counter <= "0000010111110110";
						WHEN "0000010111110110" =>
						DD(16, 22) <= packet_in;
						counter <= "0000010111110111";
						WHEN "0000010111110111" =>
						DD(16, 23) <= packet_in;
						counter <= "0000010111111000";
						WHEN "0000010111111000" =>
						DD(16, 24) <= packet_in;
						counter <= "0000010111111001";
						WHEN "0000010111111001" =>
						DD(16, 25) <= packet_in;
						counter <= "0000010111111010";
						WHEN "0000010111111010" =>
						DD(16, 26) <= packet_in;
						counter <= "0000010111111011";
						WHEN "0000010111111011" =>
						DD(16, 27) <= packet_in;
						counter <= "0000010111111100";
						WHEN "0000010111111100" =>
						DD(16, 28) <= packet_in;
						counter <= "0000010111111101";
						WHEN "0000010111111101" =>
						DD(16, 29) <= packet_in;
						counter <= "0000010111111110";
						WHEN "0000010111111110" =>
						DD(16, 30) <= packet_in;
						counter <= "0000010111111111";
						WHEN "0000010111111111" =>
						DD(16, 31) <= packet_in;
						counter <= "0000011000000000";
						WHEN "0000011000000000" =>
						DD(16, 32) <= packet_in;
						counter <= "0000011000000001";
						WHEN "0000011000000001" =>
						DD(16, 33) <= packet_in;
						counter <= "0000011000000010";
						WHEN "0000011000000010" =>
						DD(16, 34) <= packet_in;
						counter <= "0000011000000011";
						WHEN "0000011000000011" =>
						DD(16, 35) <= packet_in;
						counter <= "0000011000000100";
						WHEN "0000011000000100" =>
						DD(16, 36) <= packet_in;
						counter <= "0000011000000101";
						WHEN "0000011000000101" =>
						DD(16, 37) <= packet_in;
						counter <= "0000011000000110";
						WHEN "0000011000000110" =>
						DD(16, 38) <= packet_in;
						counter <= "0000011000000111";
						WHEN "0000011000000111" =>
						DD(16, 39) <= packet_in;
						counter <= "0000011000001000";
						WHEN "0000011000001000" =>
						DD(16, 40) <= packet_in;
						counter <= "0000011000001001";
						WHEN "0000011000001001" =>
						DD(16, 41) <= packet_in;
						counter <= "0000011000001010";
						WHEN "0000011000001010" =>
						DD(16, 42) <= packet_in;
						counter <= "0000011000001011";
						WHEN "0000011000001011" =>
						DD(16, 43) <= packet_in;
						counter <= "0000011000001100";
						WHEN "0000011000001100" =>
						DD(16, 44) <= packet_in;
						counter <= "0000011000001101";
						WHEN "0000011000001101" =>
						DD(16, 45) <= packet_in;
						counter <= "0000011000001110";
						WHEN "0000011000001110" =>
						DD(16, 46) <= packet_in;
						counter <= "0000011000001111";
						WHEN "0000011000001111" =>
						DD(16, 47) <= packet_in;
						counter <= "0000011000010000";
						WHEN "0000011000010000" =>
						DD(16, 48) <= packet_in;
						counter <= "0000011000010001";
						WHEN "0000011000010001" =>
						DD(16, 49) <= packet_in;
						counter <= "0000011000010010";
						WHEN "0000011000010010" =>
						DD(16, 50) <= packet_in;
						counter <= "0000011000010011";
						WHEN "0000011000010011" =>
						DD(16, 51) <= packet_in;
						counter <= "0000011000010100";
						WHEN "0000011000010100" =>
						DD(16, 52) <= packet_in;
						counter <= "0000011000010101";
						WHEN "0000011000010101" =>
						DD(16, 53) <= packet_in;
						counter <= "0000011000010110";
						WHEN "0000011000010110" =>
						DD(16, 54) <= packet_in;
						counter <= "0000011000010111";
						WHEN "0000011000010111" =>
						DD(16, 55) <= packet_in;
						counter <= "0000011000011000";
						WHEN "0000011000011000" =>
						DD(16, 56) <= packet_in;
						counter <= "0000011000011001";
						WHEN "0000011000011001" =>
						DD(16, 57) <= packet_in;
						counter <= "0000011000011010";
						WHEN "0000011000011010" =>
						DD(16, 58) <= packet_in;
						counter <= "0000011000011011";
						WHEN "0000011000011011" =>
						DD(16, 59) <= packet_in;
						counter <= "0000011000011100";
						WHEN "0000011000011100" =>
						DD(16, 60) <= packet_in;
						counter <= "0000011000011101";
						WHEN "0000011000011101" =>
						DD(16, 61) <= packet_in;
						counter <= "0000011000011110";
						WHEN "0000011000011110" =>
						DD(16, 62) <= packet_in;
						counter <= "0000011000011111";
						WHEN "0000011000011111" =>
						DD(16, 63) <= packet_in;
						counter <= "0000011000100000";
						WHEN "0000011000100000" =>
						DD(16, 64) <= packet_in;
						counter <= "0000011000100001";
						WHEN "0000011000100001" =>
						DD(16, 65) <= packet_in;
						counter <= "0000011000100010";
						WHEN "0000011000100010" =>
						DD(16, 66) <= packet_in;
						counter <= "0000011000100011";
						WHEN "0000011000100011" =>
						DD(16, 67) <= packet_in;
						counter <= "0000011000100100";
						WHEN "0000011000100100" =>
						DD(16, 68) <= packet_in;
						counter <= "0000011000100101";
						WHEN "0000011000100101" =>
						DD(16, 69) <= packet_in;
						counter <= "0000011000100110";
						WHEN "0000011000100110" =>
						DD(16, 70) <= packet_in;
						counter <= "0000011000100111";
						WHEN "0000011000100111" =>
						DD(16, 71) <= packet_in;
						counter <= "0000011000101000";
						WHEN "0000011000101000" =>
						DD(16, 72) <= packet_in;
						counter <= "0000011000101001";
						WHEN "0000011000101001" =>
						DD(16, 73) <= packet_in;
						counter <= "0000011000101010";
						WHEN "0000011000101010" =>
						DD(16, 74) <= packet_in;
						counter <= "0000011000101011";
						WHEN "0000011000101011" =>
						DD(16, 75) <= packet_in;
						counter <= "0000011000101100";
						WHEN "0000011000101100" =>
						DD(16, 76) <= packet_in;
						counter <= "0000011000101101";
						WHEN "0000011000101101" =>
						DD(16, 77) <= packet_in;
						counter <= "0000011000101110";
						WHEN "0000011000101110" =>
						DD(16, 78) <= packet_in;
						counter <= "0000011000101111";
						WHEN "0000011000101111" =>
						DD(16, 79) <= packet_in;
						counter <= "0000011000110000";
						WHEN "0000011000110000" =>
						DD(16, 80) <= packet_in;
						counter <= "0000011000110001";
						WHEN "0000011000110001" =>
						DD(16, 81) <= packet_in;
						counter <= "0000011000110010";
						WHEN "0000011000110010" =>
						DD(16, 82) <= packet_in;
						counter <= "0000011000110011";
						WHEN "0000011000110011" =>
						DD(16, 83) <= packet_in;
						counter <= "0000011000110100";
						WHEN "0000011000110100" =>
						DD(16, 84) <= packet_in;
						counter <= "0000011000110101";
						WHEN "0000011000110101" =>
						DD(16, 85) <= packet_in;
						counter <= "0000011000110110";
						WHEN "0000011000110110" =>
						DD(16, 86) <= packet_in;
						counter <= "0000011000110111";
						WHEN "0000011000110111" =>
						DD(16, 87) <= packet_in;
						counter <= "0000011000111000";
						WHEN "0000011000111000" =>
						DD(16, 88) <= packet_in;
						counter <= "0000011000111001";
						WHEN "0000011000111001" =>
						DD(16, 89) <= packet_in;
						counter <= "0000011000111010";
						WHEN "0000011000111010" =>
						DD(16, 90) <= packet_in;
						counter <= "0000011000111011";
						WHEN "0000011000111011" =>
						DD(16, 91) <= packet_in;
						counter <= "0000011000111100";
						WHEN "0000011000111100" =>
						DD(17, 0) <= packet_in;
						counter <= "0000011000111101";
						WHEN "0000011000111101" =>
						DD(17, 1) <= packet_in;
						counter <= "0000011000111110";
						WHEN "0000011000111110" =>
						DD(17, 2) <= packet_in;
						counter <= "0000011000111111";
						WHEN "0000011000111111" =>
						DD(17, 3) <= packet_in;
						counter <= "0000011001000000";
						WHEN "0000011001000000" =>
						DD(17, 4) <= packet_in;
						counter <= "0000011001000001";
						WHEN "0000011001000001" =>
						DD(17, 5) <= packet_in;
						counter <= "0000011001000010";
						WHEN "0000011001000010" =>
						DD(17, 6) <= packet_in;
						counter <= "0000011001000011";
						WHEN "0000011001000011" =>
						DD(17, 7) <= packet_in;
						counter <= "0000011001000100";
						WHEN "0000011001000100" =>
						DD(17, 8) <= packet_in;
						counter <= "0000011001000101";
						WHEN "0000011001000101" =>
						DD(17, 9) <= packet_in;
						counter <= "0000011001000110";
						WHEN "0000011001000110" =>
						DD(17, 10) <= packet_in;
						counter <= "0000011001000111";
						WHEN "0000011001000111" =>
						DD(17, 11) <= packet_in;
						counter <= "0000011001001000";
						WHEN "0000011001001000" =>
						DD(17, 12) <= packet_in;
						counter <= "0000011001001001";
						WHEN "0000011001001001" =>
						DD(17, 13) <= packet_in;
						counter <= "0000011001001010";
						WHEN "0000011001001010" =>
						DD(17, 14) <= packet_in;
						counter <= "0000011001001011";
						WHEN "0000011001001011" =>
						DD(17, 15) <= packet_in;
						counter <= "0000011001001100";
						WHEN "0000011001001100" =>
						DD(17, 16) <= packet_in;
						counter <= "0000011001001101";
						WHEN "0000011001001101" =>
						DD(17, 17) <= packet_in;
						counter <= "0000011001001110";
						WHEN "0000011001001110" =>
						DD(17, 18) <= packet_in;
						counter <= "0000011001001111";
						WHEN "0000011001001111" =>
						DD(17, 19) <= packet_in;
						counter <= "0000011001010000";
						WHEN "0000011001010000" =>
						DD(17, 20) <= packet_in;
						counter <= "0000011001010001";
						WHEN "0000011001010001" =>
						DD(17, 21) <= packet_in;
						counter <= "0000011001010010";
						WHEN "0000011001010010" =>
						DD(17, 22) <= packet_in;
						counter <= "0000011001010011";
						WHEN "0000011001010011" =>
						DD(17, 23) <= packet_in;
						counter <= "0000011001010100";
						WHEN "0000011001010100" =>
						DD(17, 24) <= packet_in;
						counter <= "0000011001010101";
						WHEN "0000011001010101" =>
						DD(17, 25) <= packet_in;
						counter <= "0000011001010110";
						WHEN "0000011001010110" =>
						DD(17, 26) <= packet_in;
						counter <= "0000011001010111";
						WHEN "0000011001010111" =>
						DD(17, 27) <= packet_in;
						counter <= "0000011001011000";
						WHEN "0000011001011000" =>
						DD(17, 28) <= packet_in;
						counter <= "0000011001011001";
						WHEN "0000011001011001" =>
						DD(17, 29) <= packet_in;
						counter <= "0000011001011010";
						WHEN "0000011001011010" =>
						DD(17, 30) <= packet_in;
						counter <= "0000011001011011";
						WHEN "0000011001011011" =>
						DD(17, 31) <= packet_in;
						counter <= "0000011001011100";
						WHEN "0000011001011100" =>
						DD(17, 32) <= packet_in;
						counter <= "0000011001011101";
						WHEN "0000011001011101" =>
						DD(17, 33) <= packet_in;
						counter <= "0000011001011110";
						WHEN "0000011001011110" =>
						DD(17, 34) <= packet_in;
						counter <= "0000011001011111";
						WHEN "0000011001011111" =>
						DD(17, 35) <= packet_in;
						counter <= "0000011001100000";
						WHEN "0000011001100000" =>
						DD(17, 36) <= packet_in;
						counter <= "0000011001100001";
						WHEN "0000011001100001" =>
						DD(17, 37) <= packet_in;
						counter <= "0000011001100010";
						WHEN "0000011001100010" =>
						DD(17, 38) <= packet_in;
						counter <= "0000011001100011";
						WHEN "0000011001100011" =>
						DD(17, 39) <= packet_in;
						counter <= "0000011001100100";
						WHEN "0000011001100100" =>
						DD(17, 40) <= packet_in;
						counter <= "0000011001100101";
						WHEN "0000011001100101" =>
						DD(17, 41) <= packet_in;
						counter <= "0000011001100110";
						WHEN "0000011001100110" =>
						DD(17, 42) <= packet_in;
						counter <= "0000011001100111";
						WHEN "0000011001100111" =>
						DD(17, 43) <= packet_in;
						counter <= "0000011001101000";
						WHEN "0000011001101000" =>
						DD(17, 44) <= packet_in;
						counter <= "0000011001101001";
						WHEN "0000011001101001" =>
						DD(17, 45) <= packet_in;
						counter <= "0000011001101010";
						WHEN "0000011001101010" =>
						DD(17, 46) <= packet_in;
						counter <= "0000011001101011";
						WHEN "0000011001101011" =>
						DD(17, 47) <= packet_in;
						counter <= "0000011001101100";
						WHEN "0000011001101100" =>
						DD(17, 48) <= packet_in;
						counter <= "0000011001101101";
						WHEN "0000011001101101" =>
						DD(17, 49) <= packet_in;
						counter <= "0000011001101110";
						WHEN "0000011001101110" =>
						DD(17, 50) <= packet_in;
						counter <= "0000011001101111";
						WHEN "0000011001101111" =>
						DD(17, 51) <= packet_in;
						counter <= "0000011001110000";
						WHEN "0000011001110000" =>
						DD(17, 52) <= packet_in;
						counter <= "0000011001110001";
						WHEN "0000011001110001" =>
						DD(17, 53) <= packet_in;
						counter <= "0000011001110010";
						WHEN "0000011001110010" =>
						DD(17, 54) <= packet_in;
						counter <= "0000011001110011";
						WHEN "0000011001110011" =>
						DD(17, 55) <= packet_in;
						counter <= "0000011001110100";
						WHEN "0000011001110100" =>
						DD(17, 56) <= packet_in;
						counter <= "0000011001110101";
						WHEN "0000011001110101" =>
						DD(17, 57) <= packet_in;
						counter <= "0000011001110110";
						WHEN "0000011001110110" =>
						DD(17, 58) <= packet_in;
						counter <= "0000011001110111";
						WHEN "0000011001110111" =>
						DD(17, 59) <= packet_in;
						counter <= "0000011001111000";
						WHEN "0000011001111000" =>
						DD(17, 60) <= packet_in;
						counter <= "0000011001111001";
						WHEN "0000011001111001" =>
						DD(17, 61) <= packet_in;
						counter <= "0000011001111010";
						WHEN "0000011001111010" =>
						DD(17, 62) <= packet_in;
						counter <= "0000011001111011";
						WHEN "0000011001111011" =>
						DD(17, 63) <= packet_in;
						counter <= "0000011001111100";
						WHEN "0000011001111100" =>
						DD(17, 64) <= packet_in;
						counter <= "0000011001111101";
						WHEN "0000011001111101" =>
						DD(17, 65) <= packet_in;
						counter <= "0000011001111110";
						WHEN "0000011001111110" =>
						DD(17, 66) <= packet_in;
						counter <= "0000011001111111";
						WHEN "0000011001111111" =>
						DD(17, 67) <= packet_in;
						counter <= "0000011010000000";
						WHEN "0000011010000000" =>
						DD(17, 68) <= packet_in;
						counter <= "0000011010000001";
						WHEN "0000011010000001" =>
						DD(17, 69) <= packet_in;
						counter <= "0000011010000010";
						WHEN "0000011010000010" =>
						DD(17, 70) <= packet_in;
						counter <= "0000011010000011";
						WHEN "0000011010000011" =>
						DD(17, 71) <= packet_in;
						counter <= "0000011010000100";
						WHEN "0000011010000100" =>
						DD(17, 72) <= packet_in;
						counter <= "0000011010000101";
						WHEN "0000011010000101" =>
						DD(17, 73) <= packet_in;
						counter <= "0000011010000110";
						WHEN "0000011010000110" =>
						DD(17, 74) <= packet_in;
						counter <= "0000011010000111";
						WHEN "0000011010000111" =>
						DD(17, 75) <= packet_in;
						counter <= "0000011010001000";
						WHEN "0000011010001000" =>
						DD(17, 76) <= packet_in;
						counter <= "0000011010001001";
						WHEN "0000011010001001" =>
						DD(17, 77) <= packet_in;
						counter <= "0000011010001010";
						WHEN "0000011010001010" =>
						DD(17, 78) <= packet_in;
						counter <= "0000011010001011";
						WHEN "0000011010001011" =>
						DD(17, 79) <= packet_in;
						counter <= "0000011010001100";
						WHEN "0000011010001100" =>
						DD(17, 80) <= packet_in;
						counter <= "0000011010001101";
						WHEN "0000011010001101" =>
						DD(17, 81) <= packet_in;
						counter <= "0000011010001110";
						WHEN "0000011010001110" =>
						DD(17, 82) <= packet_in;
						counter <= "0000011010001111";
						WHEN "0000011010001111" =>
						DD(17, 83) <= packet_in;
						counter <= "0000011010010000";
						WHEN "0000011010010000" =>
						DD(17, 84) <= packet_in;
						counter <= "0000011010010001";
						WHEN "0000011010010001" =>
						DD(17, 85) <= packet_in;
						counter <= "0000011010010010";
						WHEN "0000011010010010" =>
						DD(17, 86) <= packet_in;
						counter <= "0000011010010011";
						WHEN "0000011010010011" =>
						DD(17, 87) <= packet_in;
						counter <= "0000011010010100";
						WHEN "0000011010010100" =>
						DD(17, 88) <= packet_in;
						counter <= "0000011010010101";
						WHEN "0000011010010101" =>
						DD(17, 89) <= packet_in;
						counter <= "0000011010010110";
						WHEN "0000011010010110" =>
						DD(17, 90) <= packet_in;
						counter <= "0000011010010111";
						WHEN "0000011010010111" =>
						DD(17, 91) <= packet_in;
						counter <= "0000011010011000";
						WHEN "0000011010011000" =>
						DD(18, 0) <= packet_in;
						counter <= "0000011010011001";
						WHEN "0000011010011001" =>
						DD(18, 1) <= packet_in;
						counter <= "0000011010011010";
						WHEN "0000011010011010" =>
						DD(18, 2) <= packet_in;
						counter <= "0000011010011011";
						WHEN "0000011010011011" =>
						DD(18, 3) <= packet_in;
						counter <= "0000011010011100";
						WHEN "0000011010011100" =>
						DD(18, 4) <= packet_in;
						counter <= "0000011010011101";
						WHEN "0000011010011101" =>
						DD(18, 5) <= packet_in;
						counter <= "0000011010011110";
						WHEN "0000011010011110" =>
						DD(18, 6) <= packet_in;
						counter <= "0000011010011111";
						WHEN "0000011010011111" =>
						DD(18, 7) <= packet_in;
						counter <= "0000011010100000";
						WHEN "0000011010100000" =>
						DD(18, 8) <= packet_in;
						counter <= "0000011010100001";
						WHEN "0000011010100001" =>
						DD(18, 9) <= packet_in;
						counter <= "0000011010100010";
						WHEN "0000011010100010" =>
						DD(18, 10) <= packet_in;
						counter <= "0000011010100011";
						WHEN "0000011010100011" =>
						DD(18, 11) <= packet_in;
						counter <= "0000011010100100";
						WHEN "0000011010100100" =>
						DD(18, 12) <= packet_in;
						counter <= "0000011010100101";
						WHEN "0000011010100101" =>
						DD(18, 13) <= packet_in;
						counter <= "0000011010100110";
						WHEN "0000011010100110" =>
						DD(18, 14) <= packet_in;
						counter <= "0000011010100111";
						WHEN "0000011010100111" =>
						DD(18, 15) <= packet_in;
						counter <= "0000011010101000";
						WHEN "0000011010101000" =>
						DD(18, 16) <= packet_in;
						counter <= "0000011010101001";
						WHEN "0000011010101001" =>
						DD(18, 17) <= packet_in;
						counter <= "0000011010101010";
						WHEN "0000011010101010" =>
						DD(18, 18) <= packet_in;
						counter <= "0000011010101011";
						WHEN "0000011010101011" =>
						DD(18, 19) <= packet_in;
						counter <= "0000011010101100";
						WHEN "0000011010101100" =>
						DD(18, 20) <= packet_in;
						counter <= "0000011010101101";
						WHEN "0000011010101101" =>
						DD(18, 21) <= packet_in;
						counter <= "0000011010101110";
						WHEN "0000011010101110" =>
						DD(18, 22) <= packet_in;
						counter <= "0000011010101111";
						WHEN "0000011010101111" =>
						DD(18, 23) <= packet_in;
						counter <= "0000011010110000";
						WHEN "0000011010110000" =>
						DD(18, 24) <= packet_in;
						counter <= "0000011010110001";
						WHEN "0000011010110001" =>
						DD(18, 25) <= packet_in;
						counter <= "0000011010110010";
						WHEN "0000011010110010" =>
						DD(18, 26) <= packet_in;
						counter <= "0000011010110011";
						WHEN "0000011010110011" =>
						DD(18, 27) <= packet_in;
						counter <= "0000011010110100";
						WHEN "0000011010110100" =>
						DD(18, 28) <= packet_in;
						counter <= "0000011010110101";
						WHEN "0000011010110101" =>
						DD(18, 29) <= packet_in;
						counter <= "0000011010110110";
						WHEN "0000011010110110" =>
						DD(18, 30) <= packet_in;
						counter <= "0000011010110111";
						WHEN "0000011010110111" =>
						DD(18, 31) <= packet_in;
						counter <= "0000011010111000";
						WHEN "0000011010111000" =>
						DD(18, 32) <= packet_in;
						counter <= "0000011010111001";
						WHEN "0000011010111001" =>
						DD(18, 33) <= packet_in;
						counter <= "0000011010111010";
						WHEN "0000011010111010" =>
						DD(18, 34) <= packet_in;
						counter <= "0000011010111011";
						WHEN "0000011010111011" =>
						DD(18, 35) <= packet_in;
						counter <= "0000011010111100";
						WHEN "0000011010111100" =>
						DD(18, 36) <= packet_in;
						counter <= "0000011010111101";
						WHEN "0000011010111101" =>
						DD(18, 37) <= packet_in;
						counter <= "0000011010111110";
						WHEN "0000011010111110" =>
						DD(18, 38) <= packet_in;
						counter <= "0000011010111111";
						WHEN "0000011010111111" =>
						DD(18, 39) <= packet_in;
						counter <= "0000011011000000";
						WHEN "0000011011000000" =>
						DD(18, 40) <= packet_in;
						counter <= "0000011011000001";
						WHEN "0000011011000001" =>
						DD(18, 41) <= packet_in;
						counter <= "0000011011000010";
						WHEN "0000011011000010" =>
						DD(18, 42) <= packet_in;
						counter <= "0000011011000011";
						WHEN "0000011011000011" =>
						DD(18, 43) <= packet_in;
						counter <= "0000011011000100";
						WHEN "0000011011000100" =>
						DD(18, 44) <= packet_in;
						counter <= "0000011011000101";
						WHEN "0000011011000101" =>
						DD(18, 45) <= packet_in;
						counter <= "0000011011000110";
						WHEN "0000011011000110" =>
						DD(18, 46) <= packet_in;
						counter <= "0000011011000111";
						WHEN "0000011011000111" =>
						DD(18, 47) <= packet_in;
						counter <= "0000011011001000";
						WHEN "0000011011001000" =>
						DD(18, 48) <= packet_in;
						counter <= "0000011011001001";
						WHEN "0000011011001001" =>
						DD(18, 49) <= packet_in;
						counter <= "0000011011001010";
						WHEN "0000011011001010" =>
						DD(18, 50) <= packet_in;
						counter <= "0000011011001011";
						WHEN "0000011011001011" =>
						DD(18, 51) <= packet_in;
						counter <= "0000011011001100";
						WHEN "0000011011001100" =>
						DD(18, 52) <= packet_in;
						counter <= "0000011011001101";
						WHEN "0000011011001101" =>
						DD(18, 53) <= packet_in;
						counter <= "0000011011001110";
						WHEN "0000011011001110" =>
						DD(18, 54) <= packet_in;
						counter <= "0000011011001111";
						WHEN "0000011011001111" =>
						DD(18, 55) <= packet_in;
						counter <= "0000011011010000";
						WHEN "0000011011010000" =>
						DD(18, 56) <= packet_in;
						counter <= "0000011011010001";
						WHEN "0000011011010001" =>
						DD(18, 57) <= packet_in;
						counter <= "0000011011010010";
						WHEN "0000011011010010" =>
						DD(18, 58) <= packet_in;
						counter <= "0000011011010011";
						WHEN "0000011011010011" =>
						DD(18, 59) <= packet_in;
						counter <= "0000011011010100";
						WHEN "0000011011010100" =>
						DD(18, 60) <= packet_in;
						counter <= "0000011011010101";
						WHEN "0000011011010101" =>
						DD(18, 61) <= packet_in;
						counter <= "0000011011010110";
						WHEN "0000011011010110" =>
						DD(18, 62) <= packet_in;
						counter <= "0000011011010111";
						WHEN "0000011011010111" =>
						DD(18, 63) <= packet_in;
						counter <= "0000011011011000";
						WHEN "0000011011011000" =>
						DD(18, 64) <= packet_in;
						counter <= "0000011011011001";
						WHEN "0000011011011001" =>
						DD(18, 65) <= packet_in;
						counter <= "0000011011011010";
						WHEN "0000011011011010" =>
						DD(18, 66) <= packet_in;
						counter <= "0000011011011011";
						WHEN "0000011011011011" =>
						DD(18, 67) <= packet_in;
						counter <= "0000011011011100";
						WHEN "0000011011011100" =>
						DD(18, 68) <= packet_in;
						counter <= "0000011011011101";
						WHEN "0000011011011101" =>
						DD(18, 69) <= packet_in;
						counter <= "0000011011011110";
						WHEN "0000011011011110" =>
						DD(18, 70) <= packet_in;
						counter <= "0000011011011111";
						WHEN "0000011011011111" =>
						DD(18, 71) <= packet_in;
						counter <= "0000011011100000";
						WHEN "0000011011100000" =>
						DD(18, 72) <= packet_in;
						counter <= "0000011011100001";
						WHEN "0000011011100001" =>
						DD(18, 73) <= packet_in;
						counter <= "0000011011100010";
						WHEN "0000011011100010" =>
						DD(18, 74) <= packet_in;
						counter <= "0000011011100011";
						WHEN "0000011011100011" =>
						DD(18, 75) <= packet_in;
						counter <= "0000011011100100";
						WHEN "0000011011100100" =>
						DD(18, 76) <= packet_in;
						counter <= "0000011011100101";
						WHEN "0000011011100101" =>
						DD(18, 77) <= packet_in;
						counter <= "0000011011100110";
						WHEN "0000011011100110" =>
						DD(18, 78) <= packet_in;
						counter <= "0000011011100111";
						WHEN "0000011011100111" =>
						DD(18, 79) <= packet_in;
						counter <= "0000011011101000";
						WHEN "0000011011101000" =>
						DD(18, 80) <= packet_in;
						counter <= "0000011011101001";
						WHEN "0000011011101001" =>
						DD(18, 81) <= packet_in;
						counter <= "0000011011101010";
						WHEN "0000011011101010" =>
						DD(18, 82) <= packet_in;
						counter <= "0000011011101011";
						WHEN "0000011011101011" =>
						DD(18, 83) <= packet_in;
						counter <= "0000011011101100";
						WHEN "0000011011101100" =>
						DD(18, 84) <= packet_in;
						counter <= "0000011011101101";
						WHEN "0000011011101101" =>
						DD(18, 85) <= packet_in;
						counter <= "0000011011101110";
						WHEN "0000011011101110" =>
						DD(18, 86) <= packet_in;
						counter <= "0000011011101111";
						WHEN "0000011011101111" =>
						DD(18, 87) <= packet_in;
						counter <= "0000011011110000";
						WHEN "0000011011110000" =>
						DD(18, 88) <= packet_in;
						counter <= "0000011011110001";
						WHEN "0000011011110001" =>
						DD(18, 89) <= packet_in;
						counter <= "0000011011110010";
						WHEN "0000011011110010" =>
						DD(18, 90) <= packet_in;
						counter <= "0000011011110011";
						WHEN "0000011011110011" =>
						DD(18, 91) <= packet_in;
						counter <= "0000011011110100";
						WHEN "0000011011110100" =>
						DD(19, 0) <= packet_in;
						counter <= "0000011011110101";
						WHEN "0000011011110101" =>
						DD(19, 1) <= packet_in;
						counter <= "0000011011110110";
						WHEN "0000011011110110" =>
						DD(19, 2) <= packet_in;
						counter <= "0000011011110111";
						WHEN "0000011011110111" =>
						DD(19, 3) <= packet_in;
						counter <= "0000011011111000";
						WHEN "0000011011111000" =>
						DD(19, 4) <= packet_in;
						counter <= "0000011011111001";
						WHEN "0000011011111001" =>
						DD(19, 5) <= packet_in;
						counter <= "0000011011111010";
						WHEN "0000011011111010" =>
						DD(19, 6) <= packet_in;
						counter <= "0000011011111011";
						WHEN "0000011011111011" =>
						DD(19, 7) <= packet_in;
						counter <= "0000011011111100";
						WHEN "0000011011111100" =>
						DD(19, 8) <= packet_in;
						counter <= "0000011011111101";
						WHEN "0000011011111101" =>
						DD(19, 9) <= packet_in;
						counter <= "0000011011111110";
						WHEN "0000011011111110" =>
						DD(19, 10) <= packet_in;
						counter <= "0000011011111111";
						WHEN "0000011011111111" =>
						DD(19, 11) <= packet_in;
						counter <= "0000011100000000";
						WHEN "0000011100000000" =>
						DD(19, 12) <= packet_in;
						counter <= "0000011100000001";
						WHEN "0000011100000001" =>
						DD(19, 13) <= packet_in;
						counter <= "0000011100000010";
						WHEN "0000011100000010" =>
						DD(19, 14) <= packet_in;
						counter <= "0000011100000011";
						WHEN "0000011100000011" =>
						DD(19, 15) <= packet_in;
						counter <= "0000011100000100";
						WHEN "0000011100000100" =>
						DD(19, 16) <= packet_in;
						counter <= "0000011100000101";
						WHEN "0000011100000101" =>
						DD(19, 17) <= packet_in;
						counter <= "0000011100000110";
						WHEN "0000011100000110" =>
						DD(19, 18) <= packet_in;
						counter <= "0000011100000111";
						WHEN "0000011100000111" =>
						DD(19, 19) <= packet_in;
						counter <= "0000011100001000";
						WHEN "0000011100001000" =>
						DD(19, 20) <= packet_in;
						counter <= "0000011100001001";
						WHEN "0000011100001001" =>
						DD(19, 21) <= packet_in;
						counter <= "0000011100001010";
						WHEN "0000011100001010" =>
						DD(19, 22) <= packet_in;
						counter <= "0000011100001011";
						WHEN "0000011100001011" =>
						DD(19, 23) <= packet_in;
						counter <= "0000011100001100";
						WHEN "0000011100001100" =>
						DD(19, 24) <= packet_in;
						counter <= "0000011100001101";
						WHEN "0000011100001101" =>
						DD(19, 25) <= packet_in;
						counter <= "0000011100001110";
						WHEN "0000011100001110" =>
						DD(19, 26) <= packet_in;
						counter <= "0000011100001111";
						WHEN "0000011100001111" =>
						DD(19, 27) <= packet_in;
						counter <= "0000011100010000";
						WHEN "0000011100010000" =>
						DD(19, 28) <= packet_in;
						counter <= "0000011100010001";
						WHEN "0000011100010001" =>
						DD(19, 29) <= packet_in;
						counter <= "0000011100010010";
						WHEN "0000011100010010" =>
						DD(19, 30) <= packet_in;
						counter <= "0000011100010011";
						WHEN "0000011100010011" =>
						DD(19, 31) <= packet_in;
						counter <= "0000011100010100";
						WHEN "0000011100010100" =>
						DD(19, 32) <= packet_in;
						counter <= "0000011100010101";
						WHEN "0000011100010101" =>
						DD(19, 33) <= packet_in;
						counter <= "0000011100010110";
						WHEN "0000011100010110" =>
						DD(19, 34) <= packet_in;
						counter <= "0000011100010111";
						WHEN "0000011100010111" =>
						DD(19, 35) <= packet_in;
						counter <= "0000011100011000";
						WHEN "0000011100011000" =>
						DD(19, 36) <= packet_in;
						counter <= "0000011100011001";
						WHEN "0000011100011001" =>
						DD(19, 37) <= packet_in;
						counter <= "0000011100011010";
						WHEN "0000011100011010" =>
						DD(19, 38) <= packet_in;
						counter <= "0000011100011011";
						WHEN "0000011100011011" =>
						DD(19, 39) <= packet_in;
						counter <= "0000011100011100";
						WHEN "0000011100011100" =>
						DD(19, 40) <= packet_in;
						counter <= "0000011100011101";
						WHEN "0000011100011101" =>
						DD(19, 41) <= packet_in;
						counter <= "0000011100011110";
						WHEN "0000011100011110" =>
						DD(19, 42) <= packet_in;
						counter <= "0000011100011111";
						WHEN "0000011100011111" =>
						DD(19, 43) <= packet_in;
						counter <= "0000011100100000";
						WHEN "0000011100100000" =>
						DD(19, 44) <= packet_in;
						counter <= "0000011100100001";
						WHEN "0000011100100001" =>
						DD(19, 45) <= packet_in;
						counter <= "0000011100100010";
						WHEN "0000011100100010" =>
						DD(19, 46) <= packet_in;
						counter <= "0000011100100011";
						WHEN "0000011100100011" =>
						DD(19, 47) <= packet_in;
						counter <= "0000011100100100";
						WHEN "0000011100100100" =>
						DD(19, 48) <= packet_in;
						counter <= "0000011100100101";
						WHEN "0000011100100101" =>
						DD(19, 49) <= packet_in;
						counter <= "0000011100100110";
						WHEN "0000011100100110" =>
						DD(19, 50) <= packet_in;
						counter <= "0000011100100111";
						WHEN "0000011100100111" =>
						DD(19, 51) <= packet_in;
						counter <= "0000011100101000";
						WHEN "0000011100101000" =>
						DD(19, 52) <= packet_in;
						counter <= "0000011100101001";
						WHEN "0000011100101001" =>
						DD(19, 53) <= packet_in;
						counter <= "0000011100101010";
						WHEN "0000011100101010" =>
						DD(19, 54) <= packet_in;
						counter <= "0000011100101011";
						WHEN "0000011100101011" =>
						DD(19, 55) <= packet_in;
						counter <= "0000011100101100";
						WHEN "0000011100101100" =>
						DD(19, 56) <= packet_in;
						counter <= "0000011100101101";
						WHEN "0000011100101101" =>
						DD(19, 57) <= packet_in;
						counter <= "0000011100101110";
						WHEN "0000011100101110" =>
						DD(19, 58) <= packet_in;
						counter <= "0000011100101111";
						WHEN "0000011100101111" =>
						DD(19, 59) <= packet_in;
						counter <= "0000011100110000";
						WHEN "0000011100110000" =>
						DD(19, 60) <= packet_in;
						counter <= "0000011100110001";
						WHEN "0000011100110001" =>
						DD(19, 61) <= packet_in;
						counter <= "0000011100110010";
						WHEN "0000011100110010" =>
						DD(19, 62) <= packet_in;
						counter <= "0000011100110011";
						WHEN "0000011100110011" =>
						DD(19, 63) <= packet_in;
						counter <= "0000011100110100";
						WHEN "0000011100110100" =>
						DD(19, 64) <= packet_in;
						counter <= "0000011100110101";
						WHEN "0000011100110101" =>
						DD(19, 65) <= packet_in;
						counter <= "0000011100110110";
						WHEN "0000011100110110" =>
						DD(19, 66) <= packet_in;
						counter <= "0000011100110111";
						WHEN "0000011100110111" =>
						DD(19, 67) <= packet_in;
						counter <= "0000011100111000";
						WHEN "0000011100111000" =>
						DD(19, 68) <= packet_in;
						counter <= "0000011100111001";
						WHEN "0000011100111001" =>
						DD(19, 69) <= packet_in;
						counter <= "0000011100111010";
						WHEN "0000011100111010" =>
						DD(19, 70) <= packet_in;
						counter <= "0000011100111011";
						WHEN "0000011100111011" =>
						DD(19, 71) <= packet_in;
						counter <= "0000011100111100";
						WHEN "0000011100111100" =>
						DD(19, 72) <= packet_in;
						counter <= "0000011100111101";
						WHEN "0000011100111101" =>
						DD(19, 73) <= packet_in;
						counter <= "0000011100111110";
						WHEN "0000011100111110" =>
						DD(19, 74) <= packet_in;
						counter <= "0000011100111111";
						WHEN "0000011100111111" =>
						DD(19, 75) <= packet_in;
						counter <= "0000011101000000";
						WHEN "0000011101000000" =>
						DD(19, 76) <= packet_in;
						counter <= "0000011101000001";
						WHEN "0000011101000001" =>
						DD(19, 77) <= packet_in;
						counter <= "0000011101000010";
						WHEN "0000011101000010" =>
						DD(19, 78) <= packet_in;
						counter <= "0000011101000011";
						WHEN "0000011101000011" =>
						DD(19, 79) <= packet_in;
						counter <= "0000011101000100";
						WHEN "0000011101000100" =>
						DD(19, 80) <= packet_in;
						counter <= "0000011101000101";
						WHEN "0000011101000101" =>
						DD(19, 81) <= packet_in;
						counter <= "0000011101000110";
						WHEN "0000011101000110" =>
						DD(19, 82) <= packet_in;
						counter <= "0000011101000111";
						WHEN "0000011101000111" =>
						DD(19, 83) <= packet_in;
						counter <= "0000011101001000";
						WHEN "0000011101001000" =>
						DD(19, 84) <= packet_in;
						counter <= "0000011101001001";
						WHEN "0000011101001001" =>
						DD(19, 85) <= packet_in;
						counter <= "0000011101001010";
						WHEN "0000011101001010" =>
						DD(19, 86) <= packet_in;
						counter <= "0000011101001011";
						WHEN "0000011101001011" =>
						DD(19, 87) <= packet_in;
						counter <= "0000011101001100";
						WHEN "0000011101001100" =>
						DD(19, 88) <= packet_in;
						counter <= "0000011101001101";
						WHEN "0000011101001101" =>
						DD(19, 89) <= packet_in;
						counter <= "0000011101001110";
						WHEN "0000011101001110" =>
						DD(19, 90) <= packet_in;
						counter <= "0000011101001111";
						WHEN "0000011101001111" =>
						DD(19, 91) <= packet_in;
						counter <= "0000011101010000";
						WHEN "0000011101010000" =>
						DD(20, 0) <= packet_in;
						counter <= "0000011101010001";
						WHEN "0000011101010001" =>
						DD(20, 1) <= packet_in;
						counter <= "0000011101010010";
						WHEN "0000011101010010" =>
						DD(20, 2) <= packet_in;
						counter <= "0000011101010011";
						WHEN "0000011101010011" =>
						DD(20, 3) <= packet_in;
						counter <= "0000011101010100";
						WHEN "0000011101010100" =>
						DD(20, 4) <= packet_in;
						counter <= "0000011101010101";
						WHEN "0000011101010101" =>
						DD(20, 5) <= packet_in;
						counter <= "0000011101010110";
						WHEN "0000011101010110" =>
						DD(20, 6) <= packet_in;
						counter <= "0000011101010111";
						WHEN "0000011101010111" =>
						DD(20, 7) <= packet_in;
						counter <= "0000011101011000";
						WHEN "0000011101011000" =>
						DD(20, 8) <= packet_in;
						counter <= "0000011101011001";
						WHEN "0000011101011001" =>
						DD(20, 9) <= packet_in;
						counter <= "0000011101011010";
						WHEN "0000011101011010" =>
						DD(20, 10) <= packet_in;
						counter <= "0000011101011011";
						WHEN "0000011101011011" =>
						DD(20, 11) <= packet_in;
						counter <= "0000011101011100";
						WHEN "0000011101011100" =>
						DD(20, 12) <= packet_in;
						counter <= "0000011101011101";
						WHEN "0000011101011101" =>
						DD(20, 13) <= packet_in;
						counter <= "0000011101011110";
						WHEN "0000011101011110" =>
						DD(20, 14) <= packet_in;
						counter <= "0000011101011111";
						WHEN "0000011101011111" =>
						DD(20, 15) <= packet_in;
						counter <= "0000011101100000";
						WHEN "0000011101100000" =>
						DD(20, 16) <= packet_in;
						counter <= "0000011101100001";
						WHEN "0000011101100001" =>
						DD(20, 17) <= packet_in;
						counter <= "0000011101100010";
						WHEN "0000011101100010" =>
						DD(20, 18) <= packet_in;
						counter <= "0000011101100011";
						WHEN "0000011101100011" =>
						DD(20, 19) <= packet_in;
						counter <= "0000011101100100";
						WHEN "0000011101100100" =>
						DD(20, 20) <= packet_in;
						counter <= "0000011101100101";
						WHEN "0000011101100101" =>
						DD(20, 21) <= packet_in;
						counter <= "0000011101100110";
						WHEN "0000011101100110" =>
						DD(20, 22) <= packet_in;
						counter <= "0000011101100111";
						WHEN "0000011101100111" =>
						DD(20, 23) <= packet_in;
						counter <= "0000011101101000";
						WHEN "0000011101101000" =>
						DD(20, 24) <= packet_in;
						counter <= "0000011101101001";
						WHEN "0000011101101001" =>
						DD(20, 25) <= packet_in;
						counter <= "0000011101101010";
						WHEN "0000011101101010" =>
						DD(20, 26) <= packet_in;
						counter <= "0000011101101011";
						WHEN "0000011101101011" =>
						DD(20, 27) <= packet_in;
						counter <= "0000011101101100";
						WHEN "0000011101101100" =>
						DD(20, 28) <= packet_in;
						counter <= "0000011101101101";
						WHEN "0000011101101101" =>
						DD(20, 29) <= packet_in;
						counter <= "0000011101101110";
						WHEN "0000011101101110" =>
						DD(20, 30) <= packet_in;
						counter <= "0000011101101111";
						WHEN "0000011101101111" =>
						DD(20, 31) <= packet_in;
						counter <= "0000011101110000";
						WHEN "0000011101110000" =>
						DD(20, 32) <= packet_in;
						counter <= "0000011101110001";
						WHEN "0000011101110001" =>
						DD(20, 33) <= packet_in;
						counter <= "0000011101110010";
						WHEN "0000011101110010" =>
						DD(20, 34) <= packet_in;
						counter <= "0000011101110011";
						WHEN "0000011101110011" =>
						DD(20, 35) <= packet_in;
						counter <= "0000011101110100";
						WHEN "0000011101110100" =>
						DD(20, 36) <= packet_in;
						counter <= "0000011101110101";
						WHEN "0000011101110101" =>
						DD(20, 37) <= packet_in;
						counter <= "0000011101110110";
						WHEN "0000011101110110" =>
						DD(20, 38) <= packet_in;
						counter <= "0000011101110111";
						WHEN "0000011101110111" =>
						DD(20, 39) <= packet_in;
						counter <= "0000011101111000";
						WHEN "0000011101111000" =>
						DD(20, 40) <= packet_in;
						counter <= "0000011101111001";
						WHEN "0000011101111001" =>
						DD(20, 41) <= packet_in;
						counter <= "0000011101111010";
						WHEN "0000011101111010" =>
						DD(20, 42) <= packet_in;
						counter <= "0000011101111011";
						WHEN "0000011101111011" =>
						DD(20, 43) <= packet_in;
						counter <= "0000011101111100";
						WHEN "0000011101111100" =>
						DD(20, 44) <= packet_in;
						counter <= "0000011101111101";
						WHEN "0000011101111101" =>
						DD(20, 45) <= packet_in;
						counter <= "0000011101111110";
						WHEN "0000011101111110" =>
						DD(20, 46) <= packet_in;
						counter <= "0000011101111111";
						WHEN "0000011101111111" =>
						DD(20, 47) <= packet_in;
						counter <= "0000011110000000";
						WHEN "0000011110000000" =>
						DD(20, 48) <= packet_in;
						counter <= "0000011110000001";
						WHEN "0000011110000001" =>
						DD(20, 49) <= packet_in;
						counter <= "0000011110000010";
						WHEN "0000011110000010" =>
						DD(20, 50) <= packet_in;
						counter <= "0000011110000011";
						WHEN "0000011110000011" =>
						DD(20, 51) <= packet_in;
						counter <= "0000011110000100";
						WHEN "0000011110000100" =>
						DD(20, 52) <= packet_in;
						counter <= "0000011110000101";
						WHEN "0000011110000101" =>
						DD(20, 53) <= packet_in;
						counter <= "0000011110000110";
						WHEN "0000011110000110" =>
						DD(20, 54) <= packet_in;
						counter <= "0000011110000111";
						WHEN "0000011110000111" =>
						DD(20, 55) <= packet_in;
						counter <= "0000011110001000";
						WHEN "0000011110001000" =>
						DD(20, 56) <= packet_in;
						counter <= "0000011110001001";
						WHEN "0000011110001001" =>
						DD(20, 57) <= packet_in;
						counter <= "0000011110001010";
						WHEN "0000011110001010" =>
						DD(20, 58) <= packet_in;
						counter <= "0000011110001011";
						WHEN "0000011110001011" =>
						DD(20, 59) <= packet_in;
						counter <= "0000011110001100";
						WHEN "0000011110001100" =>
						DD(20, 60) <= packet_in;
						counter <= "0000011110001101";
						WHEN "0000011110001101" =>
						DD(20, 61) <= packet_in;
						counter <= "0000011110001110";
						WHEN "0000011110001110" =>
						DD(20, 62) <= packet_in;
						counter <= "0000011110001111";
						WHEN "0000011110001111" =>
						DD(20, 63) <= packet_in;
						counter <= "0000011110010000";
						WHEN "0000011110010000" =>
						DD(20, 64) <= packet_in;
						counter <= "0000011110010001";
						WHEN "0000011110010001" =>
						DD(20, 65) <= packet_in;
						counter <= "0000011110010010";
						WHEN "0000011110010010" =>
						DD(20, 66) <= packet_in;
						counter <= "0000011110010011";
						WHEN "0000011110010011" =>
						DD(20, 67) <= packet_in;
						counter <= "0000011110010100";
						WHEN "0000011110010100" =>
						DD(20, 68) <= packet_in;
						counter <= "0000011110010101";
						WHEN "0000011110010101" =>
						DD(20, 69) <= packet_in;
						counter <= "0000011110010110";
						WHEN "0000011110010110" =>
						DD(20, 70) <= packet_in;
						counter <= "0000011110010111";
						WHEN "0000011110010111" =>
						DD(20, 71) <= packet_in;
						counter <= "0000011110011000";
						WHEN "0000011110011000" =>
						DD(20, 72) <= packet_in;
						counter <= "0000011110011001";
						WHEN "0000011110011001" =>
						DD(20, 73) <= packet_in;
						counter <= "0000011110011010";
						WHEN "0000011110011010" =>
						DD(20, 74) <= packet_in;
						counter <= "0000011110011011";
						WHEN "0000011110011011" =>
						DD(20, 75) <= packet_in;
						counter <= "0000011110011100";
						WHEN "0000011110011100" =>
						DD(20, 76) <= packet_in;
						counter <= "0000011110011101";
						WHEN "0000011110011101" =>
						DD(20, 77) <= packet_in;
						counter <= "0000011110011110";
						WHEN "0000011110011110" =>
						DD(20, 78) <= packet_in;
						counter <= "0000011110011111";
						WHEN "0000011110011111" =>
						DD(20, 79) <= packet_in;
						counter <= "0000011110100000";
						WHEN "0000011110100000" =>
						DD(20, 80) <= packet_in;
						counter <= "0000011110100001";
						WHEN "0000011110100001" =>
						DD(20, 81) <= packet_in;
						counter <= "0000011110100010";
						WHEN "0000011110100010" =>
						DD(20, 82) <= packet_in;
						counter <= "0000011110100011";
						WHEN "0000011110100011" =>
						DD(20, 83) <= packet_in;
						counter <= "0000011110100100";
						WHEN "0000011110100100" =>
						DD(20, 84) <= packet_in;
						counter <= "0000011110100101";
						WHEN "0000011110100101" =>
						DD(20, 85) <= packet_in;
						counter <= "0000011110100110";
						WHEN "0000011110100110" =>
						DD(20, 86) <= packet_in;
						counter <= "0000011110100111";
						WHEN "0000011110100111" =>
						DD(20, 87) <= packet_in;
						counter <= "0000011110101000";
						WHEN "0000011110101000" =>
						DD(20, 88) <= packet_in;
						counter <= "0000011110101001";
						WHEN "0000011110101001" =>
						DD(20, 89) <= packet_in;
						counter <= "0000011110101010";
						WHEN "0000011110101010" =>
						DD(20, 90) <= packet_in;
						counter <= "0000011110101011";
						WHEN "0000011110101011" =>
						DD(20, 91) <= packet_in;
						counter <= "0000011110101100";
						WHEN "0000011110101100" =>
						DD(21, 0) <= packet_in;
						counter <= "0000011110101101";
						WHEN "0000011110101101" =>
						DD(21, 1) <= packet_in;
						counter <= "0000011110101110";
						WHEN "0000011110101110" =>
						DD(21, 2) <= packet_in;
						counter <= "0000011110101111";
						WHEN "0000011110101111" =>
						DD(21, 3) <= packet_in;
						counter <= "0000011110110000";
						WHEN "0000011110110000" =>
						DD(21, 4) <= packet_in;
						counter <= "0000011110110001";
						WHEN "0000011110110001" =>
						DD(21, 5) <= packet_in;
						counter <= "0000011110110010";
						WHEN "0000011110110010" =>
						DD(21, 6) <= packet_in;
						counter <= "0000011110110011";
						WHEN "0000011110110011" =>
						DD(21, 7) <= packet_in;
						counter <= "0000011110110100";
						WHEN "0000011110110100" =>
						DD(21, 8) <= packet_in;
						counter <= "0000011110110101";
						WHEN "0000011110110101" =>
						DD(21, 9) <= packet_in;
						counter <= "0000011110110110";
						WHEN "0000011110110110" =>
						DD(21, 10) <= packet_in;
						counter <= "0000011110110111";
						WHEN "0000011110110111" =>
						DD(21, 11) <= packet_in;
						counter <= "0000011110111000";
						WHEN "0000011110111000" =>
						DD(21, 12) <= packet_in;
						counter <= "0000011110111001";
						WHEN "0000011110111001" =>
						DD(21, 13) <= packet_in;
						counter <= "0000011110111010";
						WHEN "0000011110111010" =>
						DD(21, 14) <= packet_in;
						counter <= "0000011110111011";
						WHEN "0000011110111011" =>
						DD(21, 15) <= packet_in;
						counter <= "0000011110111100";
						WHEN "0000011110111100" =>
						DD(21, 16) <= packet_in;
						counter <= "0000011110111101";
						WHEN "0000011110111101" =>
						DD(21, 17) <= packet_in;
						counter <= "0000011110111110";
						WHEN "0000011110111110" =>
						DD(21, 18) <= packet_in;
						counter <= "0000011110111111";
						WHEN "0000011110111111" =>
						DD(21, 19) <= packet_in;
						counter <= "0000011111000000";
						WHEN "0000011111000000" =>
						DD(21, 20) <= packet_in;
						counter <= "0000011111000001";
						WHEN "0000011111000001" =>
						DD(21, 21) <= packet_in;
						counter <= "0000011111000010";
						WHEN "0000011111000010" =>
						DD(21, 22) <= packet_in;
						counter <= "0000011111000011";
						WHEN "0000011111000011" =>
						DD(21, 23) <= packet_in;
						counter <= "0000011111000100";
						WHEN "0000011111000100" =>
						DD(21, 24) <= packet_in;
						counter <= "0000011111000101";
						WHEN "0000011111000101" =>
						DD(21, 25) <= packet_in;
						counter <= "0000011111000110";
						WHEN "0000011111000110" =>
						DD(21, 26) <= packet_in;
						counter <= "0000011111000111";
						WHEN "0000011111000111" =>
						DD(21, 27) <= packet_in;
						counter <= "0000011111001000";
						WHEN "0000011111001000" =>
						DD(21, 28) <= packet_in;
						counter <= "0000011111001001";
						WHEN "0000011111001001" =>
						DD(21, 29) <= packet_in;
						counter <= "0000011111001010";
						WHEN "0000011111001010" =>
						DD(21, 30) <= packet_in;
						counter <= "0000011111001011";
						WHEN "0000011111001011" =>
						DD(21, 31) <= packet_in;
						counter <= "0000011111001100";
						WHEN "0000011111001100" =>
						DD(21, 32) <= packet_in;
						counter <= "0000011111001101";
						WHEN "0000011111001101" =>
						DD(21, 33) <= packet_in;
						counter <= "0000011111001110";
						WHEN "0000011111001110" =>
						DD(21, 34) <= packet_in;
						counter <= "0000011111001111";
						WHEN "0000011111001111" =>
						DD(21, 35) <= packet_in;
						counter <= "0000011111010000";
						WHEN "0000011111010000" =>
						DD(21, 36) <= packet_in;
						counter <= "0000011111010001";
						WHEN "0000011111010001" =>
						DD(21, 37) <= packet_in;
						counter <= "0000011111010010";
						WHEN "0000011111010010" =>
						DD(21, 38) <= packet_in;
						counter <= "0000011111010011";
						WHEN "0000011111010011" =>
						DD(21, 39) <= packet_in;
						counter <= "0000011111010100";
						WHEN "0000011111010100" =>
						DD(21, 40) <= packet_in;
						counter <= "0000011111010101";
						WHEN "0000011111010101" =>
						DD(21, 41) <= packet_in;
						counter <= "0000011111010110";
						WHEN "0000011111010110" =>
						DD(21, 42) <= packet_in;
						counter <= "0000011111010111";
						WHEN "0000011111010111" =>
						DD(21, 43) <= packet_in;
						counter <= "0000011111011000";
						WHEN "0000011111011000" =>
						DD(21, 44) <= packet_in;
						counter <= "0000011111011001";
						WHEN "0000011111011001" =>
						DD(21, 45) <= packet_in;
						counter <= "0000011111011010";
						WHEN "0000011111011010" =>
						DD(21, 46) <= packet_in;
						counter <= "0000011111011011";
						WHEN "0000011111011011" =>
						DD(21, 47) <= packet_in;
						counter <= "0000011111011100";
						WHEN "0000011111011100" =>
						DD(21, 48) <= packet_in;
						counter <= "0000011111011101";
						WHEN "0000011111011101" =>
						DD(21, 49) <= packet_in;
						counter <= "0000011111011110";
						WHEN "0000011111011110" =>
						DD(21, 50) <= packet_in;
						counter <= "0000011111011111";
						WHEN "0000011111011111" =>
						DD(21, 51) <= packet_in;
						counter <= "0000011111100000";
						WHEN "0000011111100000" =>
						DD(21, 52) <= packet_in;
						counter <= "0000011111100001";
						WHEN "0000011111100001" =>
						DD(21, 53) <= packet_in;
						counter <= "0000011111100010";
						WHEN "0000011111100010" =>
						DD(21, 54) <= packet_in;
						counter <= "0000011111100011";
						WHEN "0000011111100011" =>
						DD(21, 55) <= packet_in;
						counter <= "0000011111100100";
						WHEN "0000011111100100" =>
						DD(21, 56) <= packet_in;
						counter <= "0000011111100101";
						WHEN "0000011111100101" =>
						DD(21, 57) <= packet_in;
						counter <= "0000011111100110";
						WHEN "0000011111100110" =>
						DD(21, 58) <= packet_in;
						counter <= "0000011111100111";
						WHEN "0000011111100111" =>
						DD(21, 59) <= packet_in;
						counter <= "0000011111101000";
						WHEN "0000011111101000" =>
						DD(21, 60) <= packet_in;
						counter <= "0000011111101001";
						WHEN "0000011111101001" =>
						DD(21, 61) <= packet_in;
						counter <= "0000011111101010";
						WHEN "0000011111101010" =>
						DD(21, 62) <= packet_in;
						counter <= "0000011111101011";
						WHEN "0000011111101011" =>
						DD(21, 63) <= packet_in;
						counter <= "0000011111101100";
						WHEN "0000011111101100" =>
						DD(21, 64) <= packet_in;
						counter <= "0000011111101101";
						WHEN "0000011111101101" =>
						DD(21, 65) <= packet_in;
						counter <= "0000011111101110";
						WHEN "0000011111101110" =>
						DD(21, 66) <= packet_in;
						counter <= "0000011111101111";
						WHEN "0000011111101111" =>
						DD(21, 67) <= packet_in;
						counter <= "0000011111110000";
						WHEN "0000011111110000" =>
						DD(21, 68) <= packet_in;
						counter <= "0000011111110001";
						WHEN "0000011111110001" =>
						DD(21, 69) <= packet_in;
						counter <= "0000011111110010";
						WHEN "0000011111110010" =>
						DD(21, 70) <= packet_in;
						counter <= "0000011111110011";
						WHEN "0000011111110011" =>
						DD(21, 71) <= packet_in;
						counter <= "0000011111110100";
						WHEN "0000011111110100" =>
						DD(21, 72) <= packet_in;
						counter <= "0000011111110101";
						WHEN "0000011111110101" =>
						DD(21, 73) <= packet_in;
						counter <= "0000011111110110";
						WHEN "0000011111110110" =>
						DD(21, 74) <= packet_in;
						counter <= "0000011111110111";
						WHEN "0000011111110111" =>
						DD(21, 75) <= packet_in;
						counter <= "0000011111111000";
						WHEN "0000011111111000" =>
						DD(21, 76) <= packet_in;
						counter <= "0000011111111001";
						WHEN "0000011111111001" =>
						DD(21, 77) <= packet_in;
						counter <= "0000011111111010";
						WHEN "0000011111111010" =>
						DD(21, 78) <= packet_in;
						counter <= "0000011111111011";
						WHEN "0000011111111011" =>
						DD(21, 79) <= packet_in;
						counter <= "0000011111111100";
						WHEN "0000011111111100" =>
						DD(21, 80) <= packet_in;
						counter <= "0000011111111101";
						WHEN "0000011111111101" =>
						DD(21, 81) <= packet_in;
						counter <= "0000011111111110";
						WHEN "0000011111111110" =>
						DD(21, 82) <= packet_in;
						counter <= "0000011111111111";
						WHEN "0000011111111111" =>
						DD(21, 83) <= packet_in;
						counter <= "0000100000000000";
						WHEN "0000100000000000" =>
						DD(21, 84) <= packet_in;
						counter <= "0000100000000001";
						WHEN "0000100000000001" =>
						DD(21, 85) <= packet_in;
						counter <= "0000100000000010";
						WHEN "0000100000000010" =>
						DD(21, 86) <= packet_in;
						counter <= "0000100000000011";
						WHEN "0000100000000011" =>
						DD(21, 87) <= packet_in;
						counter <= "0000100000000100";
						WHEN "0000100000000100" =>
						DD(21, 88) <= packet_in;
						counter <= "0000100000000101";
						WHEN "0000100000000101" =>
						DD(21, 89) <= packet_in;
						counter <= "0000100000000110";
						WHEN "0000100000000110" =>
						DD(21, 90) <= packet_in;
						counter <= "0000100000000111";
						WHEN "0000100000000111" =>
						DD(21, 91) <= packet_in;
						counter <= "0000100000001000";
						WHEN "0000100000001000" =>
						DD(22, 0) <= packet_in;
						counter <= "0000100000001001";
						WHEN "0000100000001001" =>
						DD(22, 1) <= packet_in;
						counter <= "0000100000001010";
						WHEN "0000100000001010" =>
						DD(22, 2) <= packet_in;
						counter <= "0000100000001011";
						WHEN "0000100000001011" =>
						DD(22, 3) <= packet_in;
						counter <= "0000100000001100";
						WHEN "0000100000001100" =>
						DD(22, 4) <= packet_in;
						counter <= "0000100000001101";
						WHEN "0000100000001101" =>
						DD(22, 5) <= packet_in;
						counter <= "0000100000001110";
						WHEN "0000100000001110" =>
						DD(22, 6) <= packet_in;
						counter <= "0000100000001111";
						WHEN "0000100000001111" =>
						DD(22, 7) <= packet_in;
						counter <= "0000100000010000";
						WHEN "0000100000010000" =>
						DD(22, 8) <= packet_in;
						counter <= "0000100000010001";
						WHEN "0000100000010001" =>
						DD(22, 9) <= packet_in;
						counter <= "0000100000010010";
						WHEN "0000100000010010" =>
						DD(22, 10) <= packet_in;
						counter <= "0000100000010011";
						WHEN "0000100000010011" =>
						DD(22, 11) <= packet_in;
						counter <= "0000100000010100";
						WHEN "0000100000010100" =>
						DD(22, 12) <= packet_in;
						counter <= "0000100000010101";
						WHEN "0000100000010101" =>
						DD(22, 13) <= packet_in;
						counter <= "0000100000010110";
						WHEN "0000100000010110" =>
						DD(22, 14) <= packet_in;
						counter <= "0000100000010111";
						WHEN "0000100000010111" =>
						DD(22, 15) <= packet_in;
						counter <= "0000100000011000";
						WHEN "0000100000011000" =>
						DD(22, 16) <= packet_in;
						counter <= "0000100000011001";
						WHEN "0000100000011001" =>
						DD(22, 17) <= packet_in;
						counter <= "0000100000011010";
						WHEN "0000100000011010" =>
						DD(22, 18) <= packet_in;
						counter <= "0000100000011011";
						WHEN "0000100000011011" =>
						DD(22, 19) <= packet_in;
						counter <= "0000100000011100";
						WHEN "0000100000011100" =>
						DD(22, 20) <= packet_in;
						counter <= "0000100000011101";
						WHEN "0000100000011101" =>
						DD(22, 21) <= packet_in;
						counter <= "0000100000011110";
						WHEN "0000100000011110" =>
						DD(22, 22) <= packet_in;
						counter <= "0000100000011111";
						WHEN "0000100000011111" =>
						DD(22, 23) <= packet_in;
						counter <= "0000100000100000";
						WHEN "0000100000100000" =>
						DD(22, 24) <= packet_in;
						counter <= "0000100000100001";
						WHEN "0000100000100001" =>
						DD(22, 25) <= packet_in;
						counter <= "0000100000100010";
						WHEN "0000100000100010" =>
						DD(22, 26) <= packet_in;
						counter <= "0000100000100011";
						WHEN "0000100000100011" =>
						DD(22, 27) <= packet_in;
						counter <= "0000100000100100";
						WHEN "0000100000100100" =>
						DD(22, 28) <= packet_in;
						counter <= "0000100000100101";
						WHEN "0000100000100101" =>
						DD(22, 29) <= packet_in;
						counter <= "0000100000100110";
						WHEN "0000100000100110" =>
						DD(22, 30) <= packet_in;
						counter <= "0000100000100111";
						WHEN "0000100000100111" =>
						DD(22, 31) <= packet_in;
						counter <= "0000100000101000";
						WHEN "0000100000101000" =>
						DD(22, 32) <= packet_in;
						counter <= "0000100000101001";
						WHEN "0000100000101001" =>
						DD(22, 33) <= packet_in;
						counter <= "0000100000101010";
						WHEN "0000100000101010" =>
						DD(22, 34) <= packet_in;
						counter <= "0000100000101011";
						WHEN "0000100000101011" =>
						DD(22, 35) <= packet_in;
						counter <= "0000100000101100";
						WHEN "0000100000101100" =>
						DD(22, 36) <= packet_in;
						counter <= "0000100000101101";
						WHEN "0000100000101101" =>
						DD(22, 37) <= packet_in;
						counter <= "0000100000101110";
						WHEN "0000100000101110" =>
						DD(22, 38) <= packet_in;
						counter <= "0000100000101111";
						WHEN "0000100000101111" =>
						DD(22, 39) <= packet_in;
						counter <= "0000100000110000";
						WHEN "0000100000110000" =>
						DD(22, 40) <= packet_in;
						counter <= "0000100000110001";
						WHEN "0000100000110001" =>
						DD(22, 41) <= packet_in;
						counter <= "0000100000110010";
						WHEN "0000100000110010" =>
						DD(22, 42) <= packet_in;
						counter <= "0000100000110011";
						WHEN "0000100000110011" =>
						DD(22, 43) <= packet_in;
						counter <= "0000100000110100";
						WHEN "0000100000110100" =>
						DD(22, 44) <= packet_in;
						counter <= "0000100000110101";
						WHEN "0000100000110101" =>
						DD(22, 45) <= packet_in;
						counter <= "0000100000110110";
						WHEN "0000100000110110" =>
						DD(22, 46) <= packet_in;
						counter <= "0000100000110111";
						WHEN "0000100000110111" =>
						DD(22, 47) <= packet_in;
						counter <= "0000100000111000";
						WHEN "0000100000111000" =>
						DD(22, 48) <= packet_in;
						counter <= "0000100000111001";
						WHEN "0000100000111001" =>
						DD(22, 49) <= packet_in;
						counter <= "0000100000111010";
						WHEN "0000100000111010" =>
						DD(22, 50) <= packet_in;
						counter <= "0000100000111011";
						WHEN "0000100000111011" =>
						DD(22, 51) <= packet_in;
						counter <= "0000100000111100";
						WHEN "0000100000111100" =>
						DD(22, 52) <= packet_in;
						counter <= "0000100000111101";
						WHEN "0000100000111101" =>
						DD(22, 53) <= packet_in;
						counter <= "0000100000111110";
						WHEN "0000100000111110" =>
						DD(22, 54) <= packet_in;
						counter <= "0000100000111111";
						WHEN "0000100000111111" =>
						DD(22, 55) <= packet_in;
						counter <= "0000100001000000";
						WHEN "0000100001000000" =>
						DD(22, 56) <= packet_in;
						counter <= "0000100001000001";
						WHEN "0000100001000001" =>
						DD(22, 57) <= packet_in;
						counter <= "0000100001000010";
						WHEN "0000100001000010" =>
						DD(22, 58) <= packet_in;
						counter <= "0000100001000011";
						WHEN "0000100001000011" =>
						DD(22, 59) <= packet_in;
						counter <= "0000100001000100";
						WHEN "0000100001000100" =>
						DD(22, 60) <= packet_in;
						counter <= "0000100001000101";
						WHEN "0000100001000101" =>
						DD(22, 61) <= packet_in;
						counter <= "0000100001000110";
						WHEN "0000100001000110" =>
						DD(22, 62) <= packet_in;
						counter <= "0000100001000111";
						WHEN "0000100001000111" =>
						DD(22, 63) <= packet_in;
						counter <= "0000100001001000";
						WHEN "0000100001001000" =>
						DD(22, 64) <= packet_in;
						counter <= "0000100001001001";
						WHEN "0000100001001001" =>
						DD(22, 65) <= packet_in;
						counter <= "0000100001001010";
						WHEN "0000100001001010" =>
						DD(22, 66) <= packet_in;
						counter <= "0000100001001011";
						WHEN "0000100001001011" =>
						DD(22, 67) <= packet_in;
						counter <= "0000100001001100";
						WHEN "0000100001001100" =>
						DD(22, 68) <= packet_in;
						counter <= "0000100001001101";
						WHEN "0000100001001101" =>
						DD(22, 69) <= packet_in;
						counter <= "0000100001001110";
						WHEN "0000100001001110" =>
						DD(22, 70) <= packet_in;
						counter <= "0000100001001111";
						WHEN "0000100001001111" =>
						DD(22, 71) <= packet_in;
						counter <= "0000100001010000";
						WHEN "0000100001010000" =>
						DD(22, 72) <= packet_in;
						counter <= "0000100001010001";
						WHEN "0000100001010001" =>
						DD(22, 73) <= packet_in;
						counter <= "0000100001010010";
						WHEN "0000100001010010" =>
						DD(22, 74) <= packet_in;
						counter <= "0000100001010011";
						WHEN "0000100001010011" =>
						DD(22, 75) <= packet_in;
						counter <= "0000100001010100";
						WHEN "0000100001010100" =>
						DD(22, 76) <= packet_in;
						counter <= "0000100001010101";
						WHEN "0000100001010101" =>
						DD(22, 77) <= packet_in;
						counter <= "0000100001010110";
						WHEN "0000100001010110" =>
						DD(22, 78) <= packet_in;
						counter <= "0000100001010111";
						WHEN "0000100001010111" =>
						DD(22, 79) <= packet_in;
						counter <= "0000100001011000";
						WHEN "0000100001011000" =>
						DD(22, 80) <= packet_in;
						counter <= "0000100001011001";
						WHEN "0000100001011001" =>
						DD(22, 81) <= packet_in;
						counter <= "0000100001011010";
						WHEN "0000100001011010" =>
						DD(22, 82) <= packet_in;
						counter <= "0000100001011011";
						WHEN "0000100001011011" =>
						DD(22, 83) <= packet_in;
						counter <= "0000100001011100";
						WHEN "0000100001011100" =>
						DD(22, 84) <= packet_in;
						counter <= "0000100001011101";
						WHEN "0000100001011101" =>
						DD(22, 85) <= packet_in;
						counter <= "0000100001011110";
						WHEN "0000100001011110" =>
						DD(22, 86) <= packet_in;
						counter <= "0000100001011111";
						WHEN "0000100001011111" =>
						DD(22, 87) <= packet_in;
						counter <= "0000100001100000";
						WHEN "0000100001100000" =>
						DD(22, 88) <= packet_in;
						counter <= "0000100001100001";
						WHEN "0000100001100001" =>
						DD(22, 89) <= packet_in;
						counter <= "0000100001100010";
						WHEN "0000100001100010" =>
						DD(22, 90) <= packet_in;
						counter <= "0000100001100011";
						WHEN "0000100001100011" =>
						DD(22, 91) <= packet_in;
						counter <= "0000100001100100";
						WHEN "0000100001100100" =>
						DD(23, 0) <= packet_in;
						counter <= "0000100001100101";
						WHEN "0000100001100101" =>
						DD(23, 1) <= packet_in;
						counter <= "0000100001100110";
						WHEN "0000100001100110" =>
						DD(23, 2) <= packet_in;
						counter <= "0000100001100111";
						WHEN "0000100001100111" =>
						DD(23, 3) <= packet_in;
						counter <= "0000100001101000";
						WHEN "0000100001101000" =>
						DD(23, 4) <= packet_in;
						counter <= "0000100001101001";
						WHEN "0000100001101001" =>
						DD(23, 5) <= packet_in;
						counter <= "0000100001101010";
						WHEN "0000100001101010" =>
						DD(23, 6) <= packet_in;
						counter <= "0000100001101011";
						WHEN "0000100001101011" =>
						DD(23, 7) <= packet_in;
						counter <= "0000100001101100";
						WHEN "0000100001101100" =>
						DD(23, 8) <= packet_in;
						counter <= "0000100001101101";
						WHEN "0000100001101101" =>
						DD(23, 9) <= packet_in;
						counter <= "0000100001101110";
						WHEN "0000100001101110" =>
						DD(23, 10) <= packet_in;
						counter <= "0000100001101111";
						WHEN "0000100001101111" =>
						DD(23, 11) <= packet_in;
						counter <= "0000100001110000";
						WHEN "0000100001110000" =>
						DD(23, 12) <= packet_in;
						counter <= "0000100001110001";
						WHEN "0000100001110001" =>
						DD(23, 13) <= packet_in;
						counter <= "0000100001110010";
						WHEN "0000100001110010" =>
						DD(23, 14) <= packet_in;
						counter <= "0000100001110011";
						WHEN "0000100001110011" =>
						DD(23, 15) <= packet_in;
						counter <= "0000100001110100";
						WHEN "0000100001110100" =>
						DD(23, 16) <= packet_in;
						counter <= "0000100001110101";
						WHEN "0000100001110101" =>
						DD(23, 17) <= packet_in;
						counter <= "0000100001110110";
						WHEN "0000100001110110" =>
						DD(23, 18) <= packet_in;
						counter <= "0000100001110111";
						WHEN "0000100001110111" =>
						DD(23, 19) <= packet_in;
						counter <= "0000100001111000";
						WHEN "0000100001111000" =>
						DD(23, 20) <= packet_in;
						counter <= "0000100001111001";
						WHEN "0000100001111001" =>
						DD(23, 21) <= packet_in;
						counter <= "0000100001111010";
						WHEN "0000100001111010" =>
						DD(23, 22) <= packet_in;
						counter <= "0000100001111011";
						WHEN "0000100001111011" =>
						DD(23, 23) <= packet_in;
						counter <= "0000100001111100";
						WHEN "0000100001111100" =>
						DD(23, 24) <= packet_in;
						counter <= "0000100001111101";
						WHEN "0000100001111101" =>
						DD(23, 25) <= packet_in;
						counter <= "0000100001111110";
						WHEN "0000100001111110" =>
						DD(23, 26) <= packet_in;
						counter <= "0000100001111111";
						WHEN "0000100001111111" =>
						DD(23, 27) <= packet_in;
						counter <= "0000100010000000";
						WHEN "0000100010000000" =>
						DD(23, 28) <= packet_in;
						counter <= "0000100010000001";
						WHEN "0000100010000001" =>
						DD(23, 29) <= packet_in;
						counter <= "0000100010000010";
						WHEN "0000100010000010" =>
						DD(23, 30) <= packet_in;
						counter <= "0000100010000011";
						WHEN "0000100010000011" =>
						DD(23, 31) <= packet_in;
						counter <= "0000100010000100";
						WHEN "0000100010000100" =>
						DD(23, 32) <= packet_in;
						counter <= "0000100010000101";
						WHEN "0000100010000101" =>
						DD(23, 33) <= packet_in;
						counter <= "0000100010000110";
						WHEN "0000100010000110" =>
						DD(23, 34) <= packet_in;
						counter <= "0000100010000111";
						WHEN "0000100010000111" =>
						DD(23, 35) <= packet_in;
						counter <= "0000100010001000";
						WHEN "0000100010001000" =>
						DD(23, 36) <= packet_in;
						counter <= "0000100010001001";
						WHEN "0000100010001001" =>
						DD(23, 37) <= packet_in;
						counter <= "0000100010001010";
						WHEN "0000100010001010" =>
						DD(23, 38) <= packet_in;
						counter <= "0000100010001011";
						WHEN "0000100010001011" =>
						DD(23, 39) <= packet_in;
						counter <= "0000100010001100";
						WHEN "0000100010001100" =>
						DD(23, 40) <= packet_in;
						counter <= "0000100010001101";
						WHEN "0000100010001101" =>
						DD(23, 41) <= packet_in;
						counter <= "0000100010001110";
						WHEN "0000100010001110" =>
						DD(23, 42) <= packet_in;
						counter <= "0000100010001111";
						WHEN "0000100010001111" =>
						DD(23, 43) <= packet_in;
						counter <= "0000100010010000";
						WHEN "0000100010010000" =>
						DD(23, 44) <= packet_in;
						counter <= "0000100010010001";
						WHEN "0000100010010001" =>
						DD(23, 45) <= packet_in;
						counter <= "0000100010010010";
						WHEN "0000100010010010" =>
						DD(23, 46) <= packet_in;
						counter <= "0000100010010011";
						WHEN "0000100010010011" =>
						DD(23, 47) <= packet_in;
						counter <= "0000100010010100";
						WHEN "0000100010010100" =>
						DD(23, 48) <= packet_in;
						counter <= "0000100010010101";
						WHEN "0000100010010101" =>
						DD(23, 49) <= packet_in;
						counter <= "0000100010010110";
						WHEN "0000100010010110" =>
						DD(23, 50) <= packet_in;
						counter <= "0000100010010111";
						WHEN "0000100010010111" =>
						DD(23, 51) <= packet_in;
						counter <= "0000100010011000";
						WHEN "0000100010011000" =>
						DD(23, 52) <= packet_in;
						counter <= "0000100010011001";
						WHEN "0000100010011001" =>
						DD(23, 53) <= packet_in;
						counter <= "0000100010011010";
						WHEN "0000100010011010" =>
						DD(23, 54) <= packet_in;
						counter <= "0000100010011011";
						WHEN "0000100010011011" =>
						DD(23, 55) <= packet_in;
						counter <= "0000100010011100";
						WHEN "0000100010011100" =>
						DD(23, 56) <= packet_in;
						counter <= "0000100010011101";
						WHEN "0000100010011101" =>
						DD(23, 57) <= packet_in;
						counter <= "0000100010011110";
						WHEN "0000100010011110" =>
						DD(23, 58) <= packet_in;
						counter <= "0000100010011111";
						WHEN "0000100010011111" =>
						DD(23, 59) <= packet_in;
						counter <= "0000100010100000";
						WHEN "0000100010100000" =>
						DD(23, 60) <= packet_in;
						counter <= "0000100010100001";
						WHEN "0000100010100001" =>
						DD(23, 61) <= packet_in;
						counter <= "0000100010100010";
						WHEN "0000100010100010" =>
						DD(23, 62) <= packet_in;
						counter <= "0000100010100011";
						WHEN "0000100010100011" =>
						DD(23, 63) <= packet_in;
						counter <= "0000100010100100";
						WHEN "0000100010100100" =>
						DD(23, 64) <= packet_in;
						counter <= "0000100010100101";
						WHEN "0000100010100101" =>
						DD(23, 65) <= packet_in;
						counter <= "0000100010100110";
						WHEN "0000100010100110" =>
						DD(23, 66) <= packet_in;
						counter <= "0000100010100111";
						WHEN "0000100010100111" =>
						DD(23, 67) <= packet_in;
						counter <= "0000100010101000";
						WHEN "0000100010101000" =>
						DD(23, 68) <= packet_in;
						counter <= "0000100010101001";
						WHEN "0000100010101001" =>
						DD(23, 69) <= packet_in;
						counter <= "0000100010101010";
						WHEN "0000100010101010" =>
						DD(23, 70) <= packet_in;
						counter <= "0000100010101011";
						WHEN "0000100010101011" =>
						DD(23, 71) <= packet_in;
						counter <= "0000100010101100";
						WHEN "0000100010101100" =>
						DD(23, 72) <= packet_in;
						counter <= "0000100010101101";
						WHEN "0000100010101101" =>
						DD(23, 73) <= packet_in;
						counter <= "0000100010101110";
						WHEN "0000100010101110" =>
						DD(23, 74) <= packet_in;
						counter <= "0000100010101111";
						WHEN "0000100010101111" =>
						DD(23, 75) <= packet_in;
						counter <= "0000100010110000";
						WHEN "0000100010110000" =>
						DD(23, 76) <= packet_in;
						counter <= "0000100010110001";
						WHEN "0000100010110001" =>
						DD(23, 77) <= packet_in;
						counter <= "0000100010110010";
						WHEN "0000100010110010" =>
						DD(23, 78) <= packet_in;
						counter <= "0000100010110011";
						WHEN "0000100010110011" =>
						DD(23, 79) <= packet_in;
						counter <= "0000100010110100";
						WHEN "0000100010110100" =>
						DD(23, 80) <= packet_in;
						counter <= "0000100010110101";
						WHEN "0000100010110101" =>
						DD(23, 81) <= packet_in;
						counter <= "0000100010110110";
						WHEN "0000100010110110" =>
						DD(23, 82) <= packet_in;
						counter <= "0000100010110111";
						WHEN "0000100010110111" =>
						DD(23, 83) <= packet_in;
						counter <= "0000100010111000";
						WHEN "0000100010111000" =>
						DD(23, 84) <= packet_in;
						counter <= "0000100010111001";
						WHEN "0000100010111001" =>
						DD(23, 85) <= packet_in;
						counter <= "0000100010111010";
						WHEN "0000100010111010" =>
						DD(23, 86) <= packet_in;
						counter <= "0000100010111011";
						WHEN "0000100010111011" =>
						DD(23, 87) <= packet_in;
						counter <= "0000100010111100";
						WHEN "0000100010111100" =>
						DD(23, 88) <= packet_in;
						counter <= "0000100010111101";
						WHEN "0000100010111101" =>
						DD(23, 89) <= packet_in;
						counter <= "0000100010111110";
						WHEN "0000100010111110" =>
						DD(23, 90) <= packet_in;
						counter <= "0000100010111111";
						WHEN "0000100010111111" =>
						DD(23, 91) <= packet_in;
						counter <= "0000100011000000";
						WHEN "0000100011000000" =>
						DD(24, 0) <= packet_in;
						counter <= "0000100011000001";
						WHEN "0000100011000001" =>
						DD(24, 1) <= packet_in;
						counter <= "0000100011000010";
						WHEN "0000100011000010" =>
						DD(24, 2) <= packet_in;
						counter <= "0000100011000011";
						WHEN "0000100011000011" =>
						DD(24, 3) <= packet_in;
						counter <= "0000100011000100";
						WHEN "0000100011000100" =>
						DD(24, 4) <= packet_in;
						counter <= "0000100011000101";
						WHEN "0000100011000101" =>
						DD(24, 5) <= packet_in;
						counter <= "0000100011000110";
						WHEN "0000100011000110" =>
						DD(24, 6) <= packet_in;
						counter <= "0000100011000111";
						WHEN "0000100011000111" =>
						DD(24, 7) <= packet_in;
						counter <= "0000100011001000";
						WHEN "0000100011001000" =>
						DD(24, 8) <= packet_in;
						counter <= "0000100011001001";
						WHEN "0000100011001001" =>
						DD(24, 9) <= packet_in;
						counter <= "0000100011001010";
						WHEN "0000100011001010" =>
						DD(24, 10) <= packet_in;
						counter <= "0000100011001011";
						WHEN "0000100011001011" =>
						DD(24, 11) <= packet_in;
						counter <= "0000100011001100";
						WHEN "0000100011001100" =>
						DD(24, 12) <= packet_in;
						counter <= "0000100011001101";
						WHEN "0000100011001101" =>
						DD(24, 13) <= packet_in;
						counter <= "0000100011001110";
						WHEN "0000100011001110" =>
						DD(24, 14) <= packet_in;
						counter <= "0000100011001111";
						WHEN "0000100011001111" =>
						DD(24, 15) <= packet_in;
						counter <= "0000100011010000";
						WHEN "0000100011010000" =>
						DD(24, 16) <= packet_in;
						counter <= "0000100011010001";
						WHEN "0000100011010001" =>
						DD(24, 17) <= packet_in;
						counter <= "0000100011010010";
						WHEN "0000100011010010" =>
						DD(24, 18) <= packet_in;
						counter <= "0000100011010011";
						WHEN "0000100011010011" =>
						DD(24, 19) <= packet_in;
						counter <= "0000100011010100";
						WHEN "0000100011010100" =>
						DD(24, 20) <= packet_in;
						counter <= "0000100011010101";
						WHEN "0000100011010101" =>
						DD(24, 21) <= packet_in;
						counter <= "0000100011010110";
						WHEN "0000100011010110" =>
						DD(24, 22) <= packet_in;
						counter <= "0000100011010111";
						WHEN "0000100011010111" =>
						DD(24, 23) <= packet_in;
						counter <= "0000100011011000";
						WHEN "0000100011011000" =>
						DD(24, 24) <= packet_in;
						counter <= "0000100011011001";
						WHEN "0000100011011001" =>
						DD(24, 25) <= packet_in;
						counter <= "0000100011011010";
						WHEN "0000100011011010" =>
						DD(24, 26) <= packet_in;
						counter <= "0000100011011011";
						WHEN "0000100011011011" =>
						DD(24, 27) <= packet_in;
						counter <= "0000100011011100";
						WHEN "0000100011011100" =>
						DD(24, 28) <= packet_in;
						counter <= "0000100011011101";
						WHEN "0000100011011101" =>
						DD(24, 29) <= packet_in;
						counter <= "0000100011011110";
						WHEN "0000100011011110" =>
						DD(24, 30) <= packet_in;
						counter <= "0000100011011111";
						WHEN "0000100011011111" =>
						DD(24, 31) <= packet_in;
						counter <= "0000100011100000";
						WHEN "0000100011100000" =>
						DD(24, 32) <= packet_in;
						counter <= "0000100011100001";
						WHEN "0000100011100001" =>
						DD(24, 33) <= packet_in;
						counter <= "0000100011100010";
						WHEN "0000100011100010" =>
						DD(24, 34) <= packet_in;
						counter <= "0000100011100011";
						WHEN "0000100011100011" =>
						DD(24, 35) <= packet_in;
						counter <= "0000100011100100";
						WHEN "0000100011100100" =>
						DD(24, 36) <= packet_in;
						counter <= "0000100011100101";
						WHEN "0000100011100101" =>
						DD(24, 37) <= packet_in;
						counter <= "0000100011100110";
						WHEN "0000100011100110" =>
						DD(24, 38) <= packet_in;
						counter <= "0000100011100111";
						WHEN "0000100011100111" =>
						DD(24, 39) <= packet_in;
						counter <= "0000100011101000";
						WHEN "0000100011101000" =>
						DD(24, 40) <= packet_in;
						counter <= "0000100011101001";
						WHEN "0000100011101001" =>
						DD(24, 41) <= packet_in;
						counter <= "0000100011101010";
						WHEN "0000100011101010" =>
						DD(24, 42) <= packet_in;
						counter <= "0000100011101011";
						WHEN "0000100011101011" =>
						DD(24, 43) <= packet_in;
						counter <= "0000100011101100";
						WHEN "0000100011101100" =>
						DD(24, 44) <= packet_in;
						counter <= "0000100011101101";
						WHEN "0000100011101101" =>
						DD(24, 45) <= packet_in;
						counter <= "0000100011101110";
						WHEN "0000100011101110" =>
						DD(24, 46) <= packet_in;
						counter <= "0000100011101111";
						WHEN "0000100011101111" =>
						DD(24, 47) <= packet_in;
						counter <= "0000100011110000";
						WHEN "0000100011110000" =>
						DD(24, 48) <= packet_in;
						counter <= "0000100011110001";
						WHEN "0000100011110001" =>
						DD(24, 49) <= packet_in;
						counter <= "0000100011110010";
						WHEN "0000100011110010" =>
						DD(24, 50) <= packet_in;
						counter <= "0000100011110011";
						WHEN "0000100011110011" =>
						DD(24, 51) <= packet_in;
						counter <= "0000100011110100";
						WHEN "0000100011110100" =>
						DD(24, 52) <= packet_in;
						counter <= "0000100011110101";
						WHEN "0000100011110101" =>
						DD(24, 53) <= packet_in;
						counter <= "0000100011110110";
						WHEN "0000100011110110" =>
						DD(24, 54) <= packet_in;
						counter <= "0000100011110111";
						WHEN "0000100011110111" =>
						DD(24, 55) <= packet_in;
						counter <= "0000100011111000";
						WHEN "0000100011111000" =>
						DD(24, 56) <= packet_in;
						counter <= "0000100011111001";
						WHEN "0000100011111001" =>
						DD(24, 57) <= packet_in;
						counter <= "0000100011111010";
						WHEN "0000100011111010" =>
						DD(24, 58) <= packet_in;
						counter <= "0000100011111011";
						WHEN "0000100011111011" =>
						DD(24, 59) <= packet_in;
						counter <= "0000100011111100";
						WHEN "0000100011111100" =>
						DD(24, 60) <= packet_in;
						counter <= "0000100011111101";
						WHEN "0000100011111101" =>
						DD(24, 61) <= packet_in;
						counter <= "0000100011111110";
						WHEN "0000100011111110" =>
						DD(24, 62) <= packet_in;
						counter <= "0000100011111111";
						WHEN "0000100011111111" =>
						DD(24, 63) <= packet_in;
						counter <= "0000100100000000";
						WHEN "0000100100000000" =>
						DD(24, 64) <= packet_in;
						counter <= "0000100100000001";
						WHEN "0000100100000001" =>
						DD(24, 65) <= packet_in;
						counter <= "0000100100000010";
						WHEN "0000100100000010" =>
						DD(24, 66) <= packet_in;
						counter <= "0000100100000011";
						WHEN "0000100100000011" =>
						DD(24, 67) <= packet_in;
						counter <= "0000100100000100";
						WHEN "0000100100000100" =>
						DD(24, 68) <= packet_in;
						counter <= "0000100100000101";
						WHEN "0000100100000101" =>
						DD(24, 69) <= packet_in;
						counter <= "0000100100000110";
						WHEN "0000100100000110" =>
						DD(24, 70) <= packet_in;
						counter <= "0000100100000111";
						WHEN "0000100100000111" =>
						DD(24, 71) <= packet_in;
						counter <= "0000100100001000";
						WHEN "0000100100001000" =>
						DD(24, 72) <= packet_in;
						counter <= "0000100100001001";
						WHEN "0000100100001001" =>
						DD(24, 73) <= packet_in;
						counter <= "0000100100001010";
						WHEN "0000100100001010" =>
						DD(24, 74) <= packet_in;
						counter <= "0000100100001011";
						WHEN "0000100100001011" =>
						DD(24, 75) <= packet_in;
						counter <= "0000100100001100";
						WHEN "0000100100001100" =>
						DD(24, 76) <= packet_in;
						counter <= "0000100100001101";
						WHEN "0000100100001101" =>
						DD(24, 77) <= packet_in;
						counter <= "0000100100001110";
						WHEN "0000100100001110" =>
						DD(24, 78) <= packet_in;
						counter <= "0000100100001111";
						WHEN "0000100100001111" =>
						DD(24, 79) <= packet_in;
						counter <= "0000100100010000";
						WHEN "0000100100010000" =>
						DD(24, 80) <= packet_in;
						counter <= "0000100100010001";
						WHEN "0000100100010001" =>
						DD(24, 81) <= packet_in;
						counter <= "0000100100010010";
						WHEN "0000100100010010" =>
						DD(24, 82) <= packet_in;
						counter <= "0000100100010011";
						WHEN "0000100100010011" =>
						DD(24, 83) <= packet_in;
						counter <= "0000100100010100";
						WHEN "0000100100010100" =>
						DD(24, 84) <= packet_in;
						counter <= "0000100100010101";
						WHEN "0000100100010101" =>
						DD(24, 85) <= packet_in;
						counter <= "0000100100010110";
						WHEN "0000100100010110" =>
						DD(24, 86) <= packet_in;
						counter <= "0000100100010111";
						WHEN "0000100100010111" =>
						DD(24, 87) <= packet_in;
						counter <= "0000100100011000";
						WHEN "0000100100011000" =>
						DD(24, 88) <= packet_in;
						counter <= "0000100100011001";
						WHEN "0000100100011001" =>
						DD(24, 89) <= packet_in;
						counter <= "0000100100011010";
						WHEN "0000100100011010" =>
						DD(24, 90) <= packet_in;
						counter <= "0000100100011011";
						WHEN "0000100100011011" =>
						DD(24, 91) <= packet_in;
						counter <= "0000100100011100";
						WHEN "0000100100011100" =>
						DD(25, 0) <= packet_in;
						counter <= "0000100100011101";
						WHEN "0000100100011101" =>
						DD(25, 1) <= packet_in;
						counter <= "0000100100011110";
						WHEN "0000100100011110" =>
						DD(25, 2) <= packet_in;
						counter <= "0000100100011111";
						WHEN "0000100100011111" =>
						DD(25, 3) <= packet_in;
						counter <= "0000100100100000";
						WHEN "0000100100100000" =>
						DD(25, 4) <= packet_in;
						counter <= "0000100100100001";
						WHEN "0000100100100001" =>
						DD(25, 5) <= packet_in;
						counter <= "0000100100100010";
						WHEN "0000100100100010" =>
						DD(25, 6) <= packet_in;
						counter <= "0000100100100011";
						WHEN "0000100100100011" =>
						DD(25, 7) <= packet_in;
						counter <= "0000100100100100";
						WHEN "0000100100100100" =>
						DD(25, 8) <= packet_in;
						counter <= "0000100100100101";
						WHEN "0000100100100101" =>
						DD(25, 9) <= packet_in;
						counter <= "0000100100100110";
						WHEN "0000100100100110" =>
						DD(25, 10) <= packet_in;
						counter <= "0000100100100111";
						WHEN "0000100100100111" =>
						DD(25, 11) <= packet_in;
						counter <= "0000100100101000";
						WHEN "0000100100101000" =>
						DD(25, 12) <= packet_in;
						counter <= "0000100100101001";
						WHEN "0000100100101001" =>
						DD(25, 13) <= packet_in;
						counter <= "0000100100101010";
						WHEN "0000100100101010" =>
						DD(25, 14) <= packet_in;
						counter <= "0000100100101011";
						WHEN "0000100100101011" =>
						DD(25, 15) <= packet_in;
						counter <= "0000100100101100";
						WHEN "0000100100101100" =>
						DD(25, 16) <= packet_in;
						counter <= "0000100100101101";
						WHEN "0000100100101101" =>
						DD(25, 17) <= packet_in;
						counter <= "0000100100101110";
						WHEN "0000100100101110" =>
						DD(25, 18) <= packet_in;
						counter <= "0000100100101111";
						WHEN "0000100100101111" =>
						DD(25, 19) <= packet_in;
						counter <= "0000100100110000";
						WHEN "0000100100110000" =>
						DD(25, 20) <= packet_in;
						counter <= "0000100100110001";
						WHEN "0000100100110001" =>
						DD(25, 21) <= packet_in;
						counter <= "0000100100110010";
						WHEN "0000100100110010" =>
						DD(25, 22) <= packet_in;
						counter <= "0000100100110011";
						WHEN "0000100100110011" =>
						DD(25, 23) <= packet_in;
						counter <= "0000100100110100";
						WHEN "0000100100110100" =>
						DD(25, 24) <= packet_in;
						counter <= "0000100100110101";
						WHEN "0000100100110101" =>
						DD(25, 25) <= packet_in;
						counter <= "0000100100110110";
						WHEN "0000100100110110" =>
						DD(25, 26) <= packet_in;
						counter <= "0000100100110111";
						WHEN "0000100100110111" =>
						DD(25, 27) <= packet_in;
						counter <= "0000100100111000";
						WHEN "0000100100111000" =>
						DD(25, 28) <= packet_in;
						counter <= "0000100100111001";
						WHEN "0000100100111001" =>
						DD(25, 29) <= packet_in;
						counter <= "0000100100111010";
						WHEN "0000100100111010" =>
						DD(25, 30) <= packet_in;
						counter <= "0000100100111011";
						WHEN "0000100100111011" =>
						DD(25, 31) <= packet_in;
						counter <= "0000100100111100";
						WHEN "0000100100111100" =>
						DD(25, 32) <= packet_in;
						counter <= "0000100100111101";
						WHEN "0000100100111101" =>
						DD(25, 33) <= packet_in;
						counter <= "0000100100111110";
						WHEN "0000100100111110" =>
						DD(25, 34) <= packet_in;
						counter <= "0000100100111111";
						WHEN "0000100100111111" =>
						DD(25, 35) <= packet_in;
						counter <= "0000100101000000";
						WHEN "0000100101000000" =>
						DD(25, 36) <= packet_in;
						counter <= "0000100101000001";
						WHEN "0000100101000001" =>
						DD(25, 37) <= packet_in;
						counter <= "0000100101000010";
						WHEN "0000100101000010" =>
						DD(25, 38) <= packet_in;
						counter <= "0000100101000011";
						WHEN "0000100101000011" =>
						DD(25, 39) <= packet_in;
						counter <= "0000100101000100";
						WHEN "0000100101000100" =>
						DD(25, 40) <= packet_in;
						counter <= "0000100101000101";
						WHEN "0000100101000101" =>
						DD(25, 41) <= packet_in;
						counter <= "0000100101000110";
						WHEN "0000100101000110" =>
						DD(25, 42) <= packet_in;
						counter <= "0000100101000111";
						WHEN "0000100101000111" =>
						DD(25, 43) <= packet_in;
						counter <= "0000100101001000";
						WHEN "0000100101001000" =>
						DD(25, 44) <= packet_in;
						counter <= "0000100101001001";
						WHEN "0000100101001001" =>
						DD(25, 45) <= packet_in;
						counter <= "0000100101001010";
						WHEN "0000100101001010" =>
						DD(25, 46) <= packet_in;
						counter <= "0000100101001011";
						WHEN "0000100101001011" =>
						DD(25, 47) <= packet_in;
						counter <= "0000100101001100";
						WHEN "0000100101001100" =>
						DD(25, 48) <= packet_in;
						counter <= "0000100101001101";
						WHEN "0000100101001101" =>
						DD(25, 49) <= packet_in;
						counter <= "0000100101001110";
						WHEN "0000100101001110" =>
						DD(25, 50) <= packet_in;
						counter <= "0000100101001111";
						WHEN "0000100101001111" =>
						DD(25, 51) <= packet_in;
						counter <= "0000100101010000";
						WHEN "0000100101010000" =>
						DD(25, 52) <= packet_in;
						counter <= "0000100101010001";
						WHEN "0000100101010001" =>
						DD(25, 53) <= packet_in;
						counter <= "0000100101010010";
						WHEN "0000100101010010" =>
						DD(25, 54) <= packet_in;
						counter <= "0000100101010011";
						WHEN "0000100101010011" =>
						DD(25, 55) <= packet_in;
						counter <= "0000100101010100";
						WHEN "0000100101010100" =>
						DD(25, 56) <= packet_in;
						counter <= "0000100101010101";
						WHEN "0000100101010101" =>
						DD(25, 57) <= packet_in;
						counter <= "0000100101010110";
						WHEN "0000100101010110" =>
						DD(25, 58) <= packet_in;
						counter <= "0000100101010111";
						WHEN "0000100101010111" =>
						DD(25, 59) <= packet_in;
						counter <= "0000100101011000";
						WHEN "0000100101011000" =>
						DD(25, 60) <= packet_in;
						counter <= "0000100101011001";
						WHEN "0000100101011001" =>
						DD(25, 61) <= packet_in;
						counter <= "0000100101011010";
						WHEN "0000100101011010" =>
						DD(25, 62) <= packet_in;
						counter <= "0000100101011011";
						WHEN "0000100101011011" =>
						DD(25, 63) <= packet_in;
						counter <= "0000100101011100";
						WHEN "0000100101011100" =>
						DD(25, 64) <= packet_in;
						counter <= "0000100101011101";
						WHEN "0000100101011101" =>
						DD(25, 65) <= packet_in;
						counter <= "0000100101011110";
						WHEN "0000100101011110" =>
						DD(25, 66) <= packet_in;
						counter <= "0000100101011111";
						WHEN "0000100101011111" =>
						DD(25, 67) <= packet_in;
						counter <= "0000100101100000";
						WHEN "0000100101100000" =>
						DD(25, 68) <= packet_in;
						counter <= "0000100101100001";
						WHEN "0000100101100001" =>
						DD(25, 69) <= packet_in;
						counter <= "0000100101100010";
						WHEN "0000100101100010" =>
						DD(25, 70) <= packet_in;
						counter <= "0000100101100011";
						WHEN "0000100101100011" =>
						DD(25, 71) <= packet_in;
						counter <= "0000100101100100";
						WHEN "0000100101100100" =>
						DD(25, 72) <= packet_in;
						counter <= "0000100101100101";
						WHEN "0000100101100101" =>
						DD(25, 73) <= packet_in;
						counter <= "0000100101100110";
						WHEN "0000100101100110" =>
						DD(25, 74) <= packet_in;
						counter <= "0000100101100111";
						WHEN "0000100101100111" =>
						DD(25, 75) <= packet_in;
						counter <= "0000100101101000";
						WHEN "0000100101101000" =>
						DD(25, 76) <= packet_in;
						counter <= "0000100101101001";
						WHEN "0000100101101001" =>
						DD(25, 77) <= packet_in;
						counter <= "0000100101101010";
						WHEN "0000100101101010" =>
						DD(25, 78) <= packet_in;
						counter <= "0000100101101011";
						WHEN "0000100101101011" =>
						DD(25, 79) <= packet_in;
						counter <= "0000100101101100";
						WHEN "0000100101101100" =>
						DD(25, 80) <= packet_in;
						counter <= "0000100101101101";
						WHEN "0000100101101101" =>
						DD(25, 81) <= packet_in;
						counter <= "0000100101101110";
						WHEN "0000100101101110" =>
						DD(25, 82) <= packet_in;
						counter <= "0000100101101111";
						WHEN "0000100101101111" =>
						DD(25, 83) <= packet_in;
						counter <= "0000100101110000";
						WHEN "0000100101110000" =>
						DD(25, 84) <= packet_in;
						counter <= "0000100101110001";
						WHEN "0000100101110001" =>
						DD(25, 85) <= packet_in;
						counter <= "0000100101110010";
						WHEN "0000100101110010" =>
						DD(25, 86) <= packet_in;
						counter <= "0000100101110011";
						WHEN "0000100101110011" =>
						DD(25, 87) <= packet_in;
						counter <= "0000100101110100";
						WHEN "0000100101110100" =>
						DD(25, 88) <= packet_in;
						counter <= "0000100101110101";
						WHEN "0000100101110101" =>
						DD(25, 89) <= packet_in;
						counter <= "0000100101110110";
						WHEN "0000100101110110" =>
						DD(25, 90) <= packet_in;
						counter <= "0000100101110111";
						WHEN "0000100101110111" =>
						DD(25, 91) <= packet_in;
						counter <= "0000100101111000";
						WHEN "0000100101111000" =>
						DD(26, 0) <= packet_in;
						counter <= "0000100101111001";
						WHEN "0000100101111001" =>
						DD(26, 1) <= packet_in;
						counter <= "0000100101111010";
						WHEN "0000100101111010" =>
						DD(26, 2) <= packet_in;
						counter <= "0000100101111011";
						WHEN "0000100101111011" =>
						DD(26, 3) <= packet_in;
						counter <= "0000100101111100";
						WHEN "0000100101111100" =>
						DD(26, 4) <= packet_in;
						counter <= "0000100101111101";
						WHEN "0000100101111101" =>
						DD(26, 5) <= packet_in;
						counter <= "0000100101111110";
						WHEN "0000100101111110" =>
						DD(26, 6) <= packet_in;
						counter <= "0000100101111111";
						WHEN "0000100101111111" =>
						DD(26, 7) <= packet_in;
						counter <= "0000100110000000";
						WHEN "0000100110000000" =>
						DD(26, 8) <= packet_in;
						counter <= "0000100110000001";
						WHEN "0000100110000001" =>
						DD(26, 9) <= packet_in;
						counter <= "0000100110000010";
						WHEN "0000100110000010" =>
						DD(26, 10) <= packet_in;
						counter <= "0000100110000011";
						WHEN "0000100110000011" =>
						DD(26, 11) <= packet_in;
						counter <= "0000100110000100";
						WHEN "0000100110000100" =>
						DD(26, 12) <= packet_in;
						counter <= "0000100110000101";
						WHEN "0000100110000101" =>
						DD(26, 13) <= packet_in;
						counter <= "0000100110000110";
						WHEN "0000100110000110" =>
						DD(26, 14) <= packet_in;
						counter <= "0000100110000111";
						WHEN "0000100110000111" =>
						DD(26, 15) <= packet_in;
						counter <= "0000100110001000";
						WHEN "0000100110001000" =>
						DD(26, 16) <= packet_in;
						counter <= "0000100110001001";
						WHEN "0000100110001001" =>
						DD(26, 17) <= packet_in;
						counter <= "0000100110001010";
						WHEN "0000100110001010" =>
						DD(26, 18) <= packet_in;
						counter <= "0000100110001011";
						WHEN "0000100110001011" =>
						DD(26, 19) <= packet_in;
						counter <= "0000100110001100";
						WHEN "0000100110001100" =>
						DD(26, 20) <= packet_in;
						counter <= "0000100110001101";
						WHEN "0000100110001101" =>
						DD(26, 21) <= packet_in;
						counter <= "0000100110001110";
						WHEN "0000100110001110" =>
						DD(26, 22) <= packet_in;
						counter <= "0000100110001111";
						WHEN "0000100110001111" =>
						DD(26, 23) <= packet_in;
						counter <= "0000100110010000";
						WHEN "0000100110010000" =>
						DD(26, 24) <= packet_in;
						counter <= "0000100110010001";
						WHEN "0000100110010001" =>
						DD(26, 25) <= packet_in;
						counter <= "0000100110010010";
						WHEN "0000100110010010" =>
						DD(26, 26) <= packet_in;
						counter <= "0000100110010011";
						WHEN "0000100110010011" =>
						DD(26, 27) <= packet_in;
						counter <= "0000100110010100";
						WHEN "0000100110010100" =>
						DD(26, 28) <= packet_in;
						counter <= "0000100110010101";
						WHEN "0000100110010101" =>
						DD(26, 29) <= packet_in;
						counter <= "0000100110010110";
						WHEN "0000100110010110" =>
						DD(26, 30) <= packet_in;
						counter <= "0000100110010111";
						WHEN "0000100110010111" =>
						DD(26, 31) <= packet_in;
						counter <= "0000100110011000";
						WHEN "0000100110011000" =>
						DD(26, 32) <= packet_in;
						counter <= "0000100110011001";
						WHEN "0000100110011001" =>
						DD(26, 33) <= packet_in;
						counter <= "0000100110011010";
						WHEN "0000100110011010" =>
						DD(26, 34) <= packet_in;
						counter <= "0000100110011011";
						WHEN "0000100110011011" =>
						DD(26, 35) <= packet_in;
						counter <= "0000100110011100";
						WHEN "0000100110011100" =>
						DD(26, 36) <= packet_in;
						counter <= "0000100110011101";
						WHEN "0000100110011101" =>
						DD(26, 37) <= packet_in;
						counter <= "0000100110011110";
						WHEN "0000100110011110" =>
						DD(26, 38) <= packet_in;
						counter <= "0000100110011111";
						WHEN "0000100110011111" =>
						DD(26, 39) <= packet_in;
						counter <= "0000100110100000";
						WHEN "0000100110100000" =>
						DD(26, 40) <= packet_in;
						counter <= "0000100110100001";
						WHEN "0000100110100001" =>
						DD(26, 41) <= packet_in;
						counter <= "0000100110100010";
						WHEN "0000100110100010" =>
						DD(26, 42) <= packet_in;
						counter <= "0000100110100011";
						WHEN "0000100110100011" =>
						DD(26, 43) <= packet_in;
						counter <= "0000100110100100";
						WHEN "0000100110100100" =>
						DD(26, 44) <= packet_in;
						counter <= "0000100110100101";
						WHEN "0000100110100101" =>
						DD(26, 45) <= packet_in;
						counter <= "0000100110100110";
						WHEN "0000100110100110" =>
						DD(26, 46) <= packet_in;
						counter <= "0000100110100111";
						WHEN "0000100110100111" =>
						DD(26, 47) <= packet_in;
						counter <= "0000100110101000";
						WHEN "0000100110101000" =>
						DD(26, 48) <= packet_in;
						counter <= "0000100110101001";
						WHEN "0000100110101001" =>
						DD(26, 49) <= packet_in;
						counter <= "0000100110101010";
						WHEN "0000100110101010" =>
						DD(26, 50) <= packet_in;
						counter <= "0000100110101011";
						WHEN "0000100110101011" =>
						DD(26, 51) <= packet_in;
						counter <= "0000100110101100";
						WHEN "0000100110101100" =>
						DD(26, 52) <= packet_in;
						counter <= "0000100110101101";
						WHEN "0000100110101101" =>
						DD(26, 53) <= packet_in;
						counter <= "0000100110101110";
						WHEN "0000100110101110" =>
						DD(26, 54) <= packet_in;
						counter <= "0000100110101111";
						WHEN "0000100110101111" =>
						DD(26, 55) <= packet_in;
						counter <= "0000100110110000";
						WHEN "0000100110110000" =>
						DD(26, 56) <= packet_in;
						counter <= "0000100110110001";
						WHEN "0000100110110001" =>
						DD(26, 57) <= packet_in;
						counter <= "0000100110110010";
						WHEN "0000100110110010" =>
						DD(26, 58) <= packet_in;
						counter <= "0000100110110011";
						WHEN "0000100110110011" =>
						DD(26, 59) <= packet_in;
						counter <= "0000100110110100";
						WHEN "0000100110110100" =>
						DD(26, 60) <= packet_in;
						counter <= "0000100110110101";
						WHEN "0000100110110101" =>
						DD(26, 61) <= packet_in;
						counter <= "0000100110110110";
						WHEN "0000100110110110" =>
						DD(26, 62) <= packet_in;
						counter <= "0000100110110111";
						WHEN "0000100110110111" =>
						DD(26, 63) <= packet_in;
						counter <= "0000100110111000";
						WHEN "0000100110111000" =>
						DD(26, 64) <= packet_in;
						counter <= "0000100110111001";
						WHEN "0000100110111001" =>
						DD(26, 65) <= packet_in;
						counter <= "0000100110111010";
						WHEN "0000100110111010" =>
						DD(26, 66) <= packet_in;
						counter <= "0000100110111011";
						WHEN "0000100110111011" =>
						DD(26, 67) <= packet_in;
						counter <= "0000100110111100";
						WHEN "0000100110111100" =>
						DD(26, 68) <= packet_in;
						counter <= "0000100110111101";
						WHEN "0000100110111101" =>
						DD(26, 69) <= packet_in;
						counter <= "0000100110111110";
						WHEN "0000100110111110" =>
						DD(26, 70) <= packet_in;
						counter <= "0000100110111111";
						WHEN "0000100110111111" =>
						DD(26, 71) <= packet_in;
						counter <= "0000100111000000";
						WHEN "0000100111000000" =>
						DD(26, 72) <= packet_in;
						counter <= "0000100111000001";
						WHEN "0000100111000001" =>
						DD(26, 73) <= packet_in;
						counter <= "0000100111000010";
						WHEN "0000100111000010" =>
						DD(26, 74) <= packet_in;
						counter <= "0000100111000011";
						WHEN "0000100111000011" =>
						DD(26, 75) <= packet_in;
						counter <= "0000100111000100";
						WHEN "0000100111000100" =>
						DD(26, 76) <= packet_in;
						counter <= "0000100111000101";
						WHEN "0000100111000101" =>
						DD(26, 77) <= packet_in;
						counter <= "0000100111000110";
						WHEN "0000100111000110" =>
						DD(26, 78) <= packet_in;
						counter <= "0000100111000111";
						WHEN "0000100111000111" =>
						DD(26, 79) <= packet_in;
						counter <= "0000100111001000";
						WHEN "0000100111001000" =>
						DD(26, 80) <= packet_in;
						counter <= "0000100111001001";
						WHEN "0000100111001001" =>
						DD(26, 81) <= packet_in;
						counter <= "0000100111001010";
						WHEN "0000100111001010" =>
						DD(26, 82) <= packet_in;
						counter <= "0000100111001011";
						WHEN "0000100111001011" =>
						DD(26, 83) <= packet_in;
						counter <= "0000100111001100";
						WHEN "0000100111001100" =>
						DD(26, 84) <= packet_in;
						counter <= "0000100111001101";
						WHEN "0000100111001101" =>
						DD(26, 85) <= packet_in;
						counter <= "0000100111001110";
						WHEN "0000100111001110" =>
						DD(26, 86) <= packet_in;
						counter <= "0000100111001111";
						WHEN "0000100111001111" =>
						DD(26, 87) <= packet_in;
						counter <= "0000100111010000";
						WHEN "0000100111010000" =>
						DD(26, 88) <= packet_in;
						counter <= "0000100111010001";
						WHEN "0000100111010001" =>
						DD(26, 89) <= packet_in;
						counter <= "0000100111010010";
						WHEN "0000100111010010" =>
						DD(26, 90) <= packet_in;
						counter <= "0000100111010011";
						WHEN "0000100111010011" =>
						DD(26, 91) <= packet_in;
						counter <= "0000100111010100";
						WHEN "0000100111010100" =>
						DD(27, 0) <= packet_in;
						counter <= "0000100111010101";
						WHEN "0000100111010101" =>
						DD(27, 1) <= packet_in;
						counter <= "0000100111010110";
						WHEN "0000100111010110" =>
						DD(27, 2) <= packet_in;
						counter <= "0000100111010111";
						WHEN "0000100111010111" =>
						DD(27, 3) <= packet_in;
						counter <= "0000100111011000";
						WHEN "0000100111011000" =>
						DD(27, 4) <= packet_in;
						counter <= "0000100111011001";
						WHEN "0000100111011001" =>
						DD(27, 5) <= packet_in;
						counter <= "0000100111011010";
						WHEN "0000100111011010" =>
						DD(27, 6) <= packet_in;
						counter <= "0000100111011011";
						WHEN "0000100111011011" =>
						DD(27, 7) <= packet_in;
						counter <= "0000100111011100";
						WHEN "0000100111011100" =>
						DD(27, 8) <= packet_in;
						counter <= "0000100111011101";
						WHEN "0000100111011101" =>
						DD(27, 9) <= packet_in;
						counter <= "0000100111011110";
						WHEN "0000100111011110" =>
						DD(27, 10) <= packet_in;
						counter <= "0000100111011111";
						WHEN "0000100111011111" =>
						DD(27, 11) <= packet_in;
						counter <= "0000100111100000";
						WHEN "0000100111100000" =>
						DD(27, 12) <= packet_in;
						counter <= "0000100111100001";
						WHEN "0000100111100001" =>
						DD(27, 13) <= packet_in;
						counter <= "0000100111100010";
						WHEN "0000100111100010" =>
						DD(27, 14) <= packet_in;
						counter <= "0000100111100011";
						WHEN "0000100111100011" =>
						DD(27, 15) <= packet_in;
						counter <= "0000100111100100";
						WHEN "0000100111100100" =>
						DD(27, 16) <= packet_in;
						counter <= "0000100111100101";
						WHEN "0000100111100101" =>
						DD(27, 17) <= packet_in;
						counter <= "0000100111100110";
						WHEN "0000100111100110" =>
						DD(27, 18) <= packet_in;
						counter <= "0000100111100111";
						WHEN "0000100111100111" =>
						DD(27, 19) <= packet_in;
						counter <= "0000100111101000";
						WHEN "0000100111101000" =>
						DD(27, 20) <= packet_in;
						counter <= "0000100111101001";
						WHEN "0000100111101001" =>
						DD(27, 21) <= packet_in;
						counter <= "0000100111101010";
						WHEN "0000100111101010" =>
						DD(27, 22) <= packet_in;
						counter <= "0000100111101011";
						WHEN "0000100111101011" =>
						DD(27, 23) <= packet_in;
						counter <= "0000100111101100";
						WHEN "0000100111101100" =>
						DD(27, 24) <= packet_in;
						counter <= "0000100111101101";
						WHEN "0000100111101101" =>
						DD(27, 25) <= packet_in;
						counter <= "0000100111101110";
						WHEN "0000100111101110" =>
						DD(27, 26) <= packet_in;
						counter <= "0000100111101111";
						WHEN "0000100111101111" =>
						DD(27, 27) <= packet_in;
						counter <= "0000100111110000";
						WHEN "0000100111110000" =>
						DD(27, 28) <= packet_in;
						counter <= "0000100111110001";
						WHEN "0000100111110001" =>
						DD(27, 29) <= packet_in;
						counter <= "0000100111110010";
						WHEN "0000100111110010" =>
						DD(27, 30) <= packet_in;
						counter <= "0000100111110011";
						WHEN "0000100111110011" =>
						DD(27, 31) <= packet_in;
						counter <= "0000100111110100";
						WHEN "0000100111110100" =>
						DD(27, 32) <= packet_in;
						counter <= "0000100111110101";
						WHEN "0000100111110101" =>
						DD(27, 33) <= packet_in;
						counter <= "0000100111110110";
						WHEN "0000100111110110" =>
						DD(27, 34) <= packet_in;
						counter <= "0000100111110111";
						WHEN "0000100111110111" =>
						DD(27, 35) <= packet_in;
						counter <= "0000100111111000";
						WHEN "0000100111111000" =>
						DD(27, 36) <= packet_in;
						counter <= "0000100111111001";
						WHEN "0000100111111001" =>
						DD(27, 37) <= packet_in;
						counter <= "0000100111111010";
						WHEN "0000100111111010" =>
						DD(27, 38) <= packet_in;
						counter <= "0000100111111011";
						WHEN "0000100111111011" =>
						DD(27, 39) <= packet_in;
						counter <= "0000100111111100";
						WHEN "0000100111111100" =>
						DD(27, 40) <= packet_in;
						counter <= "0000100111111101";
						WHEN "0000100111111101" =>
						DD(27, 41) <= packet_in;
						counter <= "0000100111111110";
						WHEN "0000100111111110" =>
						DD(27, 42) <= packet_in;
						counter <= "0000100111111111";
						WHEN "0000100111111111" =>
						DD(27, 43) <= packet_in;
						counter <= "0000101000000000";
						WHEN "0000101000000000" =>
						DD(27, 44) <= packet_in;
						counter <= "0000101000000001";
						WHEN "0000101000000001" =>
						DD(27, 45) <= packet_in;
						counter <= "0000101000000010";
						WHEN "0000101000000010" =>
						DD(27, 46) <= packet_in;
						counter <= "0000101000000011";
						WHEN "0000101000000011" =>
						DD(27, 47) <= packet_in;
						counter <= "0000101000000100";
						WHEN "0000101000000100" =>
						DD(27, 48) <= packet_in;
						counter <= "0000101000000101";
						WHEN "0000101000000101" =>
						DD(27, 49) <= packet_in;
						counter <= "0000101000000110";
						WHEN "0000101000000110" =>
						DD(27, 50) <= packet_in;
						counter <= "0000101000000111";
						WHEN "0000101000000111" =>
						DD(27, 51) <= packet_in;
						counter <= "0000101000001000";
						WHEN "0000101000001000" =>
						DD(27, 52) <= packet_in;
						counter <= "0000101000001001";
						WHEN "0000101000001001" =>
						DD(27, 53) <= packet_in;
						counter <= "0000101000001010";
						WHEN "0000101000001010" =>
						DD(27, 54) <= packet_in;
						counter <= "0000101000001011";
						WHEN "0000101000001011" =>
						DD(27, 55) <= packet_in;
						counter <= "0000101000001100";
						WHEN "0000101000001100" =>
						DD(27, 56) <= packet_in;
						counter <= "0000101000001101";
						WHEN "0000101000001101" =>
						DD(27, 57) <= packet_in;
						counter <= "0000101000001110";
						WHEN "0000101000001110" =>
						DD(27, 58) <= packet_in;
						counter <= "0000101000001111";
						WHEN "0000101000001111" =>
						DD(27, 59) <= packet_in;
						counter <= "0000101000010000";
						WHEN "0000101000010000" =>
						DD(27, 60) <= packet_in;
						counter <= "0000101000010001";
						WHEN "0000101000010001" =>
						DD(27, 61) <= packet_in;
						counter <= "0000101000010010";
						WHEN "0000101000010010" =>
						DD(27, 62) <= packet_in;
						counter <= "0000101000010011";
						WHEN "0000101000010011" =>
						DD(27, 63) <= packet_in;
						counter <= "0000101000010100";
						WHEN "0000101000010100" =>
						DD(27, 64) <= packet_in;
						counter <= "0000101000010101";
						WHEN "0000101000010101" =>
						DD(27, 65) <= packet_in;
						counter <= "0000101000010110";
						WHEN "0000101000010110" =>
						DD(27, 66) <= packet_in;
						counter <= "0000101000010111";
						WHEN "0000101000010111" =>
						DD(27, 67) <= packet_in;
						counter <= "0000101000011000";
						WHEN "0000101000011000" =>
						DD(27, 68) <= packet_in;
						counter <= "0000101000011001";
						WHEN "0000101000011001" =>
						DD(27, 69) <= packet_in;
						counter <= "0000101000011010";
						WHEN "0000101000011010" =>
						DD(27, 70) <= packet_in;
						counter <= "0000101000011011";
						WHEN "0000101000011011" =>
						DD(27, 71) <= packet_in;
						counter <= "0000101000011100";
						WHEN "0000101000011100" =>
						DD(27, 72) <= packet_in;
						counter <= "0000101000011101";
						WHEN "0000101000011101" =>
						DD(27, 73) <= packet_in;
						counter <= "0000101000011110";
						WHEN "0000101000011110" =>
						DD(27, 74) <= packet_in;
						counter <= "0000101000011111";
						WHEN "0000101000011111" =>
						DD(27, 75) <= packet_in;
						counter <= "0000101000100000";
						WHEN "0000101000100000" =>
						DD(27, 76) <= packet_in;
						counter <= "0000101000100001";
						WHEN "0000101000100001" =>
						DD(27, 77) <= packet_in;
						counter <= "0000101000100010";
						WHEN "0000101000100010" =>
						DD(27, 78) <= packet_in;
						counter <= "0000101000100011";
						WHEN "0000101000100011" =>
						DD(27, 79) <= packet_in;
						counter <= "0000101000100100";
						WHEN "0000101000100100" =>
						DD(27, 80) <= packet_in;
						counter <= "0000101000100101";
						WHEN "0000101000100101" =>
						DD(27, 81) <= packet_in;
						counter <= "0000101000100110";
						WHEN "0000101000100110" =>
						DD(27, 82) <= packet_in;
						counter <= "0000101000100111";
						WHEN "0000101000100111" =>
						DD(27, 83) <= packet_in;
						counter <= "0000101000101000";
						WHEN "0000101000101000" =>
						DD(27, 84) <= packet_in;
						counter <= "0000101000101001";
						WHEN "0000101000101001" =>
						DD(27, 85) <= packet_in;
						counter <= "0000101000101010";
						WHEN "0000101000101010" =>
						DD(27, 86) <= packet_in;
						counter <= "0000101000101011";
						WHEN "0000101000101011" =>
						DD(27, 87) <= packet_in;
						counter <= "0000101000101100";
						WHEN "0000101000101100" =>
						DD(27, 88) <= packet_in;
						counter <= "0000101000101101";
						WHEN "0000101000101101" =>
						DD(27, 89) <= packet_in;
						counter <= "0000101000101110";
						WHEN "0000101000101110" =>
						DD(27, 90) <= packet_in;
						counter <= "0000101000101111";
						WHEN "0000101000101111" =>
						DD(27, 91) <= packet_in;
						counter <= "0000101000110000";
						WHEN "0000101000110000" =>
						DD(28, 0) <= packet_in;
						counter <= "0000101000110001";
						WHEN "0000101000110001" =>
						DD(28, 1) <= packet_in;
						counter <= "0000101000110010";
						WHEN "0000101000110010" =>
						DD(28, 2) <= packet_in;
						counter <= "0000101000110011";
						WHEN "0000101000110011" =>
						DD(28, 3) <= packet_in;
						counter <= "0000101000110100";
						WHEN "0000101000110100" =>
						DD(28, 4) <= packet_in;
						counter <= "0000101000110101";
						WHEN "0000101000110101" =>
						DD(28, 5) <= packet_in;
						counter <= "0000101000110110";
						WHEN "0000101000110110" =>
						DD(28, 6) <= packet_in;
						counter <= "0000101000110111";
						WHEN "0000101000110111" =>
						DD(28, 7) <= packet_in;
						counter <= "0000101000111000";
						WHEN "0000101000111000" =>
						DD(28, 8) <= packet_in;
						counter <= "0000101000111001";
						WHEN "0000101000111001" =>
						DD(28, 9) <= packet_in;
						counter <= "0000101000111010";
						WHEN "0000101000111010" =>
						DD(28, 10) <= packet_in;
						counter <= "0000101000111011";
						WHEN "0000101000111011" =>
						DD(28, 11) <= packet_in;
						counter <= "0000101000111100";
						WHEN "0000101000111100" =>
						DD(28, 12) <= packet_in;
						counter <= "0000101000111101";
						WHEN "0000101000111101" =>
						DD(28, 13) <= packet_in;
						counter <= "0000101000111110";
						WHEN "0000101000111110" =>
						DD(28, 14) <= packet_in;
						counter <= "0000101000111111";
						WHEN "0000101000111111" =>
						DD(28, 15) <= packet_in;
						counter <= "0000101001000000";
						WHEN "0000101001000000" =>
						DD(28, 16) <= packet_in;
						counter <= "0000101001000001";
						WHEN "0000101001000001" =>
						DD(28, 17) <= packet_in;
						counter <= "0000101001000010";
						WHEN "0000101001000010" =>
						DD(28, 18) <= packet_in;
						counter <= "0000101001000011";
						WHEN "0000101001000011" =>
						DD(28, 19) <= packet_in;
						counter <= "0000101001000100";
						WHEN "0000101001000100" =>
						DD(28, 20) <= packet_in;
						counter <= "0000101001000101";
						WHEN "0000101001000101" =>
						DD(28, 21) <= packet_in;
						counter <= "0000101001000110";
						WHEN "0000101001000110" =>
						DD(28, 22) <= packet_in;
						counter <= "0000101001000111";
						WHEN "0000101001000111" =>
						DD(28, 23) <= packet_in;
						counter <= "0000101001001000";
						WHEN "0000101001001000" =>
						DD(28, 24) <= packet_in;
						counter <= "0000101001001001";
						WHEN "0000101001001001" =>
						DD(28, 25) <= packet_in;
						counter <= "0000101001001010";
						WHEN "0000101001001010" =>
						DD(28, 26) <= packet_in;
						counter <= "0000101001001011";
						WHEN "0000101001001011" =>
						DD(28, 27) <= packet_in;
						counter <= "0000101001001100";
						WHEN "0000101001001100" =>
						DD(28, 28) <= packet_in;
						counter <= "0000101001001101";
						WHEN "0000101001001101" =>
						DD(28, 29) <= packet_in;
						counter <= "0000101001001110";
						WHEN "0000101001001110" =>
						DD(28, 30) <= packet_in;
						counter <= "0000101001001111";
						WHEN "0000101001001111" =>
						DD(28, 31) <= packet_in;
						counter <= "0000101001010000";
						WHEN "0000101001010000" =>
						DD(28, 32) <= packet_in;
						counter <= "0000101001010001";
						WHEN "0000101001010001" =>
						DD(28, 33) <= packet_in;
						counter <= "0000101001010010";
						WHEN "0000101001010010" =>
						DD(28, 34) <= packet_in;
						counter <= "0000101001010011";
						WHEN "0000101001010011" =>
						DD(28, 35) <= packet_in;
						counter <= "0000101001010100";
						WHEN "0000101001010100" =>
						DD(28, 36) <= packet_in;
						counter <= "0000101001010101";
						WHEN "0000101001010101" =>
						DD(28, 37) <= packet_in;
						counter <= "0000101001010110";
						WHEN "0000101001010110" =>
						DD(28, 38) <= packet_in;
						counter <= "0000101001010111";
						WHEN "0000101001010111" =>
						DD(28, 39) <= packet_in;
						counter <= "0000101001011000";
						WHEN "0000101001011000" =>
						DD(28, 40) <= packet_in;
						counter <= "0000101001011001";
						WHEN "0000101001011001" =>
						DD(28, 41) <= packet_in;
						counter <= "0000101001011010";
						WHEN "0000101001011010" =>
						DD(28, 42) <= packet_in;
						counter <= "0000101001011011";
						WHEN "0000101001011011" =>
						DD(28, 43) <= packet_in;
						counter <= "0000101001011100";
						WHEN "0000101001011100" =>
						DD(28, 44) <= packet_in;
						counter <= "0000101001011101";
						WHEN "0000101001011101" =>
						DD(28, 45) <= packet_in;
						counter <= "0000101001011110";
						WHEN "0000101001011110" =>
						DD(28, 46) <= packet_in;
						counter <= "0000101001011111";
						WHEN "0000101001011111" =>
						DD(28, 47) <= packet_in;
						counter <= "0000101001100000";
						WHEN "0000101001100000" =>
						DD(28, 48) <= packet_in;
						counter <= "0000101001100001";
						WHEN "0000101001100001" =>
						DD(28, 49) <= packet_in;
						counter <= "0000101001100010";
						WHEN "0000101001100010" =>
						DD(28, 50) <= packet_in;
						counter <= "0000101001100011";
						WHEN "0000101001100011" =>
						DD(28, 51) <= packet_in;
						counter <= "0000101001100100";
						WHEN "0000101001100100" =>
						DD(28, 52) <= packet_in;
						counter <= "0000101001100101";
						WHEN "0000101001100101" =>
						DD(28, 53) <= packet_in;
						counter <= "0000101001100110";
						WHEN "0000101001100110" =>
						DD(28, 54) <= packet_in;
						counter <= "0000101001100111";
						WHEN "0000101001100111" =>
						DD(28, 55) <= packet_in;
						counter <= "0000101001101000";
						WHEN "0000101001101000" =>
						DD(28, 56) <= packet_in;
						counter <= "0000101001101001";
						WHEN "0000101001101001" =>
						DD(28, 57) <= packet_in;
						counter <= "0000101001101010";
						WHEN "0000101001101010" =>
						DD(28, 58) <= packet_in;
						counter <= "0000101001101011";
						WHEN "0000101001101011" =>
						DD(28, 59) <= packet_in;
						counter <= "0000101001101100";
						WHEN "0000101001101100" =>
						DD(28, 60) <= packet_in;
						counter <= "0000101001101101";
						WHEN "0000101001101101" =>
						DD(28, 61) <= packet_in;
						counter <= "0000101001101110";
						WHEN "0000101001101110" =>
						DD(28, 62) <= packet_in;
						counter <= "0000101001101111";
						WHEN "0000101001101111" =>
						DD(28, 63) <= packet_in;
						counter <= "0000101001110000";
						WHEN "0000101001110000" =>
						DD(28, 64) <= packet_in;
						counter <= "0000101001110001";
						WHEN "0000101001110001" =>
						DD(28, 65) <= packet_in;
						counter <= "0000101001110010";
						WHEN "0000101001110010" =>
						DD(28, 66) <= packet_in;
						counter <= "0000101001110011";
						WHEN "0000101001110011" =>
						DD(28, 67) <= packet_in;
						counter <= "0000101001110100";
						WHEN "0000101001110100" =>
						DD(28, 68) <= packet_in;
						counter <= "0000101001110101";
						WHEN "0000101001110101" =>
						DD(28, 69) <= packet_in;
						counter <= "0000101001110110";
						WHEN "0000101001110110" =>
						DD(28, 70) <= packet_in;
						counter <= "0000101001110111";
						WHEN "0000101001110111" =>
						DD(28, 71) <= packet_in;
						counter <= "0000101001111000";
						WHEN "0000101001111000" =>
						DD(28, 72) <= packet_in;
						counter <= "0000101001111001";
						WHEN "0000101001111001" =>
						DD(28, 73) <= packet_in;
						counter <= "0000101001111010";
						WHEN "0000101001111010" =>
						DD(28, 74) <= packet_in;
						counter <= "0000101001111011";
						WHEN "0000101001111011" =>
						DD(28, 75) <= packet_in;
						counter <= "0000101001111100";
						WHEN "0000101001111100" =>
						DD(28, 76) <= packet_in;
						counter <= "0000101001111101";
						WHEN "0000101001111101" =>
						DD(28, 77) <= packet_in;
						counter <= "0000101001111110";
						WHEN "0000101001111110" =>
						DD(28, 78) <= packet_in;
						counter <= "0000101001111111";
						WHEN "0000101001111111" =>
						DD(28, 79) <= packet_in;
						counter <= "0000101010000000";
						WHEN "0000101010000000" =>
						DD(28, 80) <= packet_in;
						counter <= "0000101010000001";
						WHEN "0000101010000001" =>
						DD(28, 81) <= packet_in;
						counter <= "0000101010000010";
						WHEN "0000101010000010" =>
						DD(28, 82) <= packet_in;
						counter <= "0000101010000011";
						WHEN "0000101010000011" =>
						DD(28, 83) <= packet_in;
						counter <= "0000101010000100";
						WHEN "0000101010000100" =>
						DD(28, 84) <= packet_in;
						counter <= "0000101010000101";
						WHEN "0000101010000101" =>
						DD(28, 85) <= packet_in;
						counter <= "0000101010000110";
						WHEN "0000101010000110" =>
						DD(28, 86) <= packet_in;
						counter <= "0000101010000111";
						WHEN "0000101010000111" =>
						DD(28, 87) <= packet_in;
						counter <= "0000101010001000";
						WHEN "0000101010001000" =>
						DD(28, 88) <= packet_in;
						counter <= "0000101010001001";
						WHEN "0000101010001001" =>
						DD(28, 89) <= packet_in;
						counter <= "0000101010001010";
						WHEN "0000101010001010" =>
						DD(28, 90) <= packet_in;
						counter <= "0000101010001011";
						WHEN "0000101010001011" =>
						DD(28, 91) <= packet_in;
						counter <= "0000101010001100";
						WHEN "0000101010001100" =>
						DD(29, 0) <= packet_in;
						counter <= "0000101010001101";
						WHEN "0000101010001101" =>
						DD(29, 1) <= packet_in;
						counter <= "0000101010001110";
						WHEN "0000101010001110" =>
						DD(29, 2) <= packet_in;
						counter <= "0000101010001111";
						WHEN "0000101010001111" =>
						DD(29, 3) <= packet_in;
						counter <= "0000101010010000";
						WHEN "0000101010010000" =>
						DD(29, 4) <= packet_in;
						counter <= "0000101010010001";
						WHEN "0000101010010001" =>
						DD(29, 5) <= packet_in;
						counter <= "0000101010010010";
						WHEN "0000101010010010" =>
						DD(29, 6) <= packet_in;
						counter <= "0000101010010011";
						WHEN "0000101010010011" =>
						DD(29, 7) <= packet_in;
						counter <= "0000101010010100";
						WHEN "0000101010010100" =>
						DD(29, 8) <= packet_in;
						counter <= "0000101010010101";
						WHEN "0000101010010101" =>
						DD(29, 9) <= packet_in;
						counter <= "0000101010010110";
						WHEN "0000101010010110" =>
						DD(29, 10) <= packet_in;
						counter <= "0000101010010111";
						WHEN "0000101010010111" =>
						DD(29, 11) <= packet_in;
						counter <= "0000101010011000";
						WHEN "0000101010011000" =>
						DD(29, 12) <= packet_in;
						counter <= "0000101010011001";
						WHEN "0000101010011001" =>
						DD(29, 13) <= packet_in;
						counter <= "0000101010011010";
						WHEN "0000101010011010" =>
						DD(29, 14) <= packet_in;
						counter <= "0000101010011011";
						WHEN "0000101010011011" =>
						DD(29, 15) <= packet_in;
						counter <= "0000101010011100";
						WHEN "0000101010011100" =>
						DD(29, 16) <= packet_in;
						counter <= "0000101010011101";
						WHEN "0000101010011101" =>
						DD(29, 17) <= packet_in;
						counter <= "0000101010011110";
						WHEN "0000101010011110" =>
						DD(29, 18) <= packet_in;
						counter <= "0000101010011111";
						WHEN "0000101010011111" =>
						DD(29, 19) <= packet_in;
						counter <= "0000101010100000";
						WHEN "0000101010100000" =>
						DD(29, 20) <= packet_in;
						counter <= "0000101010100001";
						WHEN "0000101010100001" =>
						DD(29, 21) <= packet_in;
						counter <= "0000101010100010";
						WHEN "0000101010100010" =>
						DD(29, 22) <= packet_in;
						counter <= "0000101010100011";
						WHEN "0000101010100011" =>
						DD(29, 23) <= packet_in;
						counter <= "0000101010100100";
						WHEN "0000101010100100" =>
						DD(29, 24) <= packet_in;
						counter <= "0000101010100101";
						WHEN "0000101010100101" =>
						DD(29, 25) <= packet_in;
						counter <= "0000101010100110";
						WHEN "0000101010100110" =>
						DD(29, 26) <= packet_in;
						counter <= "0000101010100111";
						WHEN "0000101010100111" =>
						DD(29, 27) <= packet_in;
						counter <= "0000101010101000";
						WHEN "0000101010101000" =>
						DD(29, 28) <= packet_in;
						counter <= "0000101010101001";
						WHEN "0000101010101001" =>
						DD(29, 29) <= packet_in;
						counter <= "0000101010101010";
						WHEN "0000101010101010" =>
						DD(29, 30) <= packet_in;
						counter <= "0000101010101011";
						WHEN "0000101010101011" =>
						DD(29, 31) <= packet_in;
						counter <= "0000101010101100";
						WHEN "0000101010101100" =>
						DD(29, 32) <= packet_in;
						counter <= "0000101010101101";
						WHEN "0000101010101101" =>
						DD(29, 33) <= packet_in;
						counter <= "0000101010101110";
						WHEN "0000101010101110" =>
						DD(29, 34) <= packet_in;
						counter <= "0000101010101111";
						WHEN "0000101010101111" =>
						DD(29, 35) <= packet_in;
						counter <= "0000101010110000";
						WHEN "0000101010110000" =>
						DD(29, 36) <= packet_in;
						counter <= "0000101010110001";
						WHEN "0000101010110001" =>
						DD(29, 37) <= packet_in;
						counter <= "0000101010110010";
						WHEN "0000101010110010" =>
						DD(29, 38) <= packet_in;
						counter <= "0000101010110011";
						WHEN "0000101010110011" =>
						DD(29, 39) <= packet_in;
						counter <= "0000101010110100";
						WHEN "0000101010110100" =>
						DD(29, 40) <= packet_in;
						counter <= "0000101010110101";
						WHEN "0000101010110101" =>
						DD(29, 41) <= packet_in;
						counter <= "0000101010110110";
						WHEN "0000101010110110" =>
						DD(29, 42) <= packet_in;
						counter <= "0000101010110111";
						WHEN "0000101010110111" =>
						DD(29, 43) <= packet_in;
						counter <= "0000101010111000";
						WHEN "0000101010111000" =>
						DD(29, 44) <= packet_in;
						counter <= "0000101010111001";
						WHEN "0000101010111001" =>
						DD(29, 45) <= packet_in;
						counter <= "0000101010111010";
						WHEN "0000101010111010" =>
						DD(29, 46) <= packet_in;
						counter <= "0000101010111011";
						WHEN "0000101010111011" =>
						DD(29, 47) <= packet_in;
						counter <= "0000101010111100";
						WHEN "0000101010111100" =>
						DD(29, 48) <= packet_in;
						counter <= "0000101010111101";
						WHEN "0000101010111101" =>
						DD(29, 49) <= packet_in;
						counter <= "0000101010111110";
						WHEN "0000101010111110" =>
						DD(29, 50) <= packet_in;
						counter <= "0000101010111111";
						WHEN "0000101010111111" =>
						DD(29, 51) <= packet_in;
						counter <= "0000101011000000";
						WHEN "0000101011000000" =>
						DD(29, 52) <= packet_in;
						counter <= "0000101011000001";
						WHEN "0000101011000001" =>
						DD(29, 53) <= packet_in;
						counter <= "0000101011000010";
						WHEN "0000101011000010" =>
						DD(29, 54) <= packet_in;
						counter <= "0000101011000011";
						WHEN "0000101011000011" =>
						DD(29, 55) <= packet_in;
						counter <= "0000101011000100";
						WHEN "0000101011000100" =>
						DD(29, 56) <= packet_in;
						counter <= "0000101011000101";
						WHEN "0000101011000101" =>
						DD(29, 57) <= packet_in;
						counter <= "0000101011000110";
						WHEN "0000101011000110" =>
						DD(29, 58) <= packet_in;
						counter <= "0000101011000111";
						WHEN "0000101011000111" =>
						DD(29, 59) <= packet_in;
						counter <= "0000101011001000";
						WHEN "0000101011001000" =>
						DD(29, 60) <= packet_in;
						counter <= "0000101011001001";
						WHEN "0000101011001001" =>
						DD(29, 61) <= packet_in;
						counter <= "0000101011001010";
						WHEN "0000101011001010" =>
						DD(29, 62) <= packet_in;
						counter <= "0000101011001011";
						WHEN "0000101011001011" =>
						DD(29, 63) <= packet_in;
						counter <= "0000101011001100";
						WHEN "0000101011001100" =>
						DD(29, 64) <= packet_in;
						counter <= "0000101011001101";
						WHEN "0000101011001101" =>
						DD(29, 65) <= packet_in;
						counter <= "0000101011001110";
						WHEN "0000101011001110" =>
						DD(29, 66) <= packet_in;
						counter <= "0000101011001111";
						WHEN "0000101011001111" =>
						DD(29, 67) <= packet_in;
						counter <= "0000101011010000";
						WHEN "0000101011010000" =>
						DD(29, 68) <= packet_in;
						counter <= "0000101011010001";
						WHEN "0000101011010001" =>
						DD(29, 69) <= packet_in;
						counter <= "0000101011010010";
						WHEN "0000101011010010" =>
						DD(29, 70) <= packet_in;
						counter <= "0000101011010011";
						WHEN "0000101011010011" =>
						DD(29, 71) <= packet_in;
						counter <= "0000101011010100";
						WHEN "0000101011010100" =>
						DD(29, 72) <= packet_in;
						counter <= "0000101011010101";
						WHEN "0000101011010101" =>
						DD(29, 73) <= packet_in;
						counter <= "0000101011010110";
						WHEN "0000101011010110" =>
						DD(29, 74) <= packet_in;
						counter <= "0000101011010111";
						WHEN "0000101011010111" =>
						DD(29, 75) <= packet_in;
						counter <= "0000101011011000";
						WHEN "0000101011011000" =>
						DD(29, 76) <= packet_in;
						counter <= "0000101011011001";
						WHEN "0000101011011001" =>
						DD(29, 77) <= packet_in;
						counter <= "0000101011011010";
						WHEN "0000101011011010" =>
						DD(29, 78) <= packet_in;
						counter <= "0000101011011011";
						WHEN "0000101011011011" =>
						DD(29, 79) <= packet_in;
						counter <= "0000101011011100";
						WHEN "0000101011011100" =>
						DD(29, 80) <= packet_in;
						counter <= "0000101011011101";
						WHEN "0000101011011101" =>
						DD(29, 81) <= packet_in;
						counter <= "0000101011011110";
						WHEN "0000101011011110" =>
						DD(29, 82) <= packet_in;
						counter <= "0000101011011111";
						WHEN "0000101011011111" =>
						DD(29, 83) <= packet_in;
						counter <= "0000101011100000";
						WHEN "0000101011100000" =>
						DD(29, 84) <= packet_in;
						counter <= "0000101011100001";
						WHEN "0000101011100001" =>
						DD(29, 85) <= packet_in;
						counter <= "0000101011100010";
						WHEN "0000101011100010" =>
						DD(29, 86) <= packet_in;
						counter <= "0000101011100011";
						WHEN "0000101011100011" =>
						DD(29, 87) <= packet_in;
						counter <= "0000101011100100";
						WHEN "0000101011100100" =>
						DD(29, 88) <= packet_in;
						counter <= "0000101011100101";
						WHEN "0000101011100101" =>
						DD(29, 89) <= packet_in;
						counter <= "0000101011100110";
						WHEN "0000101011100110" =>
						DD(29, 90) <= packet_in;
						counter <= "0000101011100111";
						WHEN "0000101011100111" =>
						DD(29, 91) <= packet_in;
						counter <= "0000101011101000";
						WHEN "0000101011101000" =>
						DD(30, 0) <= packet_in;
						counter <= "0000101011101001";
						WHEN "0000101011101001" =>
						DD(30, 1) <= packet_in;
						counter <= "0000101011101010";
						WHEN "0000101011101010" =>
						DD(30, 2) <= packet_in;
						counter <= "0000101011101011";
						WHEN "0000101011101011" =>
						DD(30, 3) <= packet_in;
						counter <= "0000101011101100";
						WHEN "0000101011101100" =>
						DD(30, 4) <= packet_in;
						counter <= "0000101011101101";
						WHEN "0000101011101101" =>
						DD(30, 5) <= packet_in;
						counter <= "0000101011101110";
						WHEN "0000101011101110" =>
						DD(30, 6) <= packet_in;
						counter <= "0000101011101111";
						WHEN "0000101011101111" =>
						DD(30, 7) <= packet_in;
						counter <= "0000101011110000";
						WHEN "0000101011110000" =>
						DD(30, 8) <= packet_in;
						counter <= "0000101011110001";
						WHEN "0000101011110001" =>
						DD(30, 9) <= packet_in;
						counter <= "0000101011110010";
						WHEN "0000101011110010" =>
						DD(30, 10) <= packet_in;
						counter <= "0000101011110011";
						WHEN "0000101011110011" =>
						DD(30, 11) <= packet_in;
						counter <= "0000101011110100";
						WHEN "0000101011110100" =>
						DD(30, 12) <= packet_in;
						counter <= "0000101011110101";
						WHEN "0000101011110101" =>
						DD(30, 13) <= packet_in;
						counter <= "0000101011110110";
						WHEN "0000101011110110" =>
						DD(30, 14) <= packet_in;
						counter <= "0000101011110111";
						WHEN "0000101011110111" =>
						DD(30, 15) <= packet_in;
						counter <= "0000101011111000";
						WHEN "0000101011111000" =>
						DD(30, 16) <= packet_in;
						counter <= "0000101011111001";
						WHEN "0000101011111001" =>
						DD(30, 17) <= packet_in;
						counter <= "0000101011111010";
						WHEN "0000101011111010" =>
						DD(30, 18) <= packet_in;
						counter <= "0000101011111011";
						WHEN "0000101011111011" =>
						DD(30, 19) <= packet_in;
						counter <= "0000101011111100";
						WHEN "0000101011111100" =>
						DD(30, 20) <= packet_in;
						counter <= "0000101011111101";
						WHEN "0000101011111101" =>
						DD(30, 21) <= packet_in;
						counter <= "0000101011111110";
						WHEN "0000101011111110" =>
						DD(30, 22) <= packet_in;
						counter <= "0000101011111111";
						WHEN "0000101011111111" =>
						DD(30, 23) <= packet_in;
						counter <= "0000101100000000";
						WHEN "0000101100000000" =>
						DD(30, 24) <= packet_in;
						counter <= "0000101100000001";
						WHEN "0000101100000001" =>
						DD(30, 25) <= packet_in;
						counter <= "0000101100000010";
						WHEN "0000101100000010" =>
						DD(30, 26) <= packet_in;
						counter <= "0000101100000011";
						WHEN "0000101100000011" =>
						DD(30, 27) <= packet_in;
						counter <= "0000101100000100";
						WHEN "0000101100000100" =>
						DD(30, 28) <= packet_in;
						counter <= "0000101100000101";
						WHEN "0000101100000101" =>
						DD(30, 29) <= packet_in;
						counter <= "0000101100000110";
						WHEN "0000101100000110" =>
						DD(30, 30) <= packet_in;
						counter <= "0000101100000111";
						WHEN "0000101100000111" =>
						DD(30, 31) <= packet_in;
						counter <= "0000101100001000";
						WHEN "0000101100001000" =>
						DD(30, 32) <= packet_in;
						counter <= "0000101100001001";
						WHEN "0000101100001001" =>
						DD(30, 33) <= packet_in;
						counter <= "0000101100001010";
						WHEN "0000101100001010" =>
						DD(30, 34) <= packet_in;
						counter <= "0000101100001011";
						WHEN "0000101100001011" =>
						DD(30, 35) <= packet_in;
						counter <= "0000101100001100";
						WHEN "0000101100001100" =>
						DD(30, 36) <= packet_in;
						counter <= "0000101100001101";
						WHEN "0000101100001101" =>
						DD(30, 37) <= packet_in;
						counter <= "0000101100001110";
						WHEN "0000101100001110" =>
						DD(30, 38) <= packet_in;
						counter <= "0000101100001111";
						WHEN "0000101100001111" =>
						DD(30, 39) <= packet_in;
						counter <= "0000101100010000";
						WHEN "0000101100010000" =>
						DD(30, 40) <= packet_in;
						counter <= "0000101100010001";
						WHEN "0000101100010001" =>
						DD(30, 41) <= packet_in;
						counter <= "0000101100010010";
						WHEN "0000101100010010" =>
						DD(30, 42) <= packet_in;
						counter <= "0000101100010011";
						WHEN "0000101100010011" =>
						DD(30, 43) <= packet_in;
						counter <= "0000101100010100";
						WHEN "0000101100010100" =>
						DD(30, 44) <= packet_in;
						counter <= "0000101100010101";
						WHEN "0000101100010101" =>
						DD(30, 45) <= packet_in;
						counter <= "0000101100010110";
						WHEN "0000101100010110" =>
						DD(30, 46) <= packet_in;
						counter <= "0000101100010111";
						WHEN "0000101100010111" =>
						DD(30, 47) <= packet_in;
						counter <= "0000101100011000";
						WHEN "0000101100011000" =>
						DD(30, 48) <= packet_in;
						counter <= "0000101100011001";
						WHEN "0000101100011001" =>
						DD(30, 49) <= packet_in;
						counter <= "0000101100011010";
						WHEN "0000101100011010" =>
						DD(30, 50) <= packet_in;
						counter <= "0000101100011011";
						WHEN "0000101100011011" =>
						DD(30, 51) <= packet_in;
						counter <= "0000101100011100";
						WHEN "0000101100011100" =>
						DD(30, 52) <= packet_in;
						counter <= "0000101100011101";
						WHEN "0000101100011101" =>
						DD(30, 53) <= packet_in;
						counter <= "0000101100011110";
						WHEN "0000101100011110" =>
						DD(30, 54) <= packet_in;
						counter <= "0000101100011111";
						WHEN "0000101100011111" =>
						DD(30, 55) <= packet_in;
						counter <= "0000101100100000";
						WHEN "0000101100100000" =>
						DD(30, 56) <= packet_in;
						counter <= "0000101100100001";
						WHEN "0000101100100001" =>
						DD(30, 57) <= packet_in;
						counter <= "0000101100100010";
						WHEN "0000101100100010" =>
						DD(30, 58) <= packet_in;
						counter <= "0000101100100011";
						WHEN "0000101100100011" =>
						DD(30, 59) <= packet_in;
						counter <= "0000101100100100";
						WHEN "0000101100100100" =>
						DD(30, 60) <= packet_in;
						counter <= "0000101100100101";
						WHEN "0000101100100101" =>
						DD(30, 61) <= packet_in;
						counter <= "0000101100100110";
						WHEN "0000101100100110" =>
						DD(30, 62) <= packet_in;
						counter <= "0000101100100111";
						WHEN "0000101100100111" =>
						DD(30, 63) <= packet_in;
						counter <= "0000101100101000";
						WHEN "0000101100101000" =>
						DD(30, 64) <= packet_in;
						counter <= "0000101100101001";
						WHEN "0000101100101001" =>
						DD(30, 65) <= packet_in;
						counter <= "0000101100101010";
						WHEN "0000101100101010" =>
						DD(30, 66) <= packet_in;
						counter <= "0000101100101011";
						WHEN "0000101100101011" =>
						DD(30, 67) <= packet_in;
						counter <= "0000101100101100";
						WHEN "0000101100101100" =>
						DD(30, 68) <= packet_in;
						counter <= "0000101100101101";
						WHEN "0000101100101101" =>
						DD(30, 69) <= packet_in;
						counter <= "0000101100101110";
						WHEN "0000101100101110" =>
						DD(30, 70) <= packet_in;
						counter <= "0000101100101111";
						WHEN "0000101100101111" =>
						DD(30, 71) <= packet_in;
						counter <= "0000101100110000";
						WHEN "0000101100110000" =>
						DD(30, 72) <= packet_in;
						counter <= "0000101100110001";
						WHEN "0000101100110001" =>
						DD(30, 73) <= packet_in;
						counter <= "0000101100110010";
						WHEN "0000101100110010" =>
						DD(30, 74) <= packet_in;
						counter <= "0000101100110011";
						WHEN "0000101100110011" =>
						DD(30, 75) <= packet_in;
						counter <= "0000101100110100";
						WHEN "0000101100110100" =>
						DD(30, 76) <= packet_in;
						counter <= "0000101100110101";
						WHEN "0000101100110101" =>
						DD(30, 77) <= packet_in;
						counter <= "0000101100110110";
						WHEN "0000101100110110" =>
						DD(30, 78) <= packet_in;
						counter <= "0000101100110111";
						WHEN "0000101100110111" =>
						DD(30, 79) <= packet_in;
						counter <= "0000101100111000";
						WHEN "0000101100111000" =>
						DD(30, 80) <= packet_in;
						counter <= "0000101100111001";
						WHEN "0000101100111001" =>
						DD(30, 81) <= packet_in;
						counter <= "0000101100111010";
						WHEN "0000101100111010" =>
						DD(30, 82) <= packet_in;
						counter <= "0000101100111011";
						WHEN "0000101100111011" =>
						DD(30, 83) <= packet_in;
						counter <= "0000101100111100";
						WHEN "0000101100111100" =>
						DD(30, 84) <= packet_in;
						counter <= "0000101100111101";
						WHEN "0000101100111101" =>
						DD(30, 85) <= packet_in;
						counter <= "0000101100111110";
						WHEN "0000101100111110" =>
						DD(30, 86) <= packet_in;
						counter <= "0000101100111111";
						WHEN "0000101100111111" =>
						DD(30, 87) <= packet_in;
						counter <= "0000101101000000";
						WHEN "0000101101000000" =>
						DD(30, 88) <= packet_in;
						counter <= "0000101101000001";
						WHEN "0000101101000001" =>
						DD(30, 89) <= packet_in;
						counter <= "0000101101000010";
						WHEN "0000101101000010" =>
						DD(30, 90) <= packet_in;
						counter <= "0000101101000011";
						WHEN "0000101101000011" =>
						DD(30, 91) <= packet_in;
						counter <= "0000101101000100";
						WHEN "0000101101000100" =>
						DD(31, 0) <= packet_in;
						counter <= "0000101101000101";
						WHEN "0000101101000101" =>
						DD(31, 1) <= packet_in;
						counter <= "0000101101000110";
						WHEN "0000101101000110" =>
						DD(31, 2) <= packet_in;
						counter <= "0000101101000111";
						WHEN "0000101101000111" =>
						DD(31, 3) <= packet_in;
						counter <= "0000101101001000";
						WHEN "0000101101001000" =>
						DD(31, 4) <= packet_in;
						counter <= "0000101101001001";
						WHEN "0000101101001001" =>
						DD(31, 5) <= packet_in;
						counter <= "0000101101001010";
						WHEN "0000101101001010" =>
						DD(31, 6) <= packet_in;
						counter <= "0000101101001011";
						WHEN "0000101101001011" =>
						DD(31, 7) <= packet_in;
						counter <= "0000101101001100";
						WHEN "0000101101001100" =>
						DD(31, 8) <= packet_in;
						counter <= "0000101101001101";
						WHEN "0000101101001101" =>
						DD(31, 9) <= packet_in;
						counter <= "0000101101001110";
						WHEN "0000101101001110" =>
						DD(31, 10) <= packet_in;
						counter <= "0000101101001111";
						WHEN "0000101101001111" =>
						DD(31, 11) <= packet_in;
						counter <= "0000101101010000";
						WHEN "0000101101010000" =>
						DD(31, 12) <= packet_in;
						counter <= "0000101101010001";
						WHEN "0000101101010001" =>
						DD(31, 13) <= packet_in;
						counter <= "0000101101010010";
						WHEN "0000101101010010" =>
						DD(31, 14) <= packet_in;
						counter <= "0000101101010011";
						WHEN "0000101101010011" =>
						DD(31, 15) <= packet_in;
						counter <= "0000101101010100";
						WHEN "0000101101010100" =>
						DD(31, 16) <= packet_in;
						counter <= "0000101101010101";
						WHEN "0000101101010101" =>
						DD(31, 17) <= packet_in;
						counter <= "0000101101010110";
						WHEN "0000101101010110" =>
						DD(31, 18) <= packet_in;
						counter <= "0000101101010111";
						WHEN "0000101101010111" =>
						DD(31, 19) <= packet_in;
						counter <= "0000101101011000";
						WHEN "0000101101011000" =>
						DD(31, 20) <= packet_in;
						counter <= "0000101101011001";
						WHEN "0000101101011001" =>
						DD(31, 21) <= packet_in;
						counter <= "0000101101011010";
						WHEN "0000101101011010" =>
						DD(31, 22) <= packet_in;
						counter <= "0000101101011011";
						WHEN "0000101101011011" =>
						DD(31, 23) <= packet_in;
						counter <= "0000101101011100";
						WHEN "0000101101011100" =>
						DD(31, 24) <= packet_in;
						counter <= "0000101101011101";
						WHEN "0000101101011101" =>
						DD(31, 25) <= packet_in;
						counter <= "0000101101011110";
						WHEN "0000101101011110" =>
						DD(31, 26) <= packet_in;
						counter <= "0000101101011111";
						WHEN "0000101101011111" =>
						DD(31, 27) <= packet_in;
						counter <= "0000101101100000";
						WHEN "0000101101100000" =>
						DD(31, 28) <= packet_in;
						counter <= "0000101101100001";
						WHEN "0000101101100001" =>
						DD(31, 29) <= packet_in;
						counter <= "0000101101100010";
						WHEN "0000101101100010" =>
						DD(31, 30) <= packet_in;
						counter <= "0000101101100011";
						WHEN "0000101101100011" =>
						DD(31, 31) <= packet_in;
						counter <= "0000101101100100";
						WHEN "0000101101100100" =>
						DD(31, 32) <= packet_in;
						counter <= "0000101101100101";
						WHEN "0000101101100101" =>
						DD(31, 33) <= packet_in;
						counter <= "0000101101100110";
						WHEN "0000101101100110" =>
						DD(31, 34) <= packet_in;
						counter <= "0000101101100111";
						WHEN "0000101101100111" =>
						DD(31, 35) <= packet_in;
						counter <= "0000101101101000";
						WHEN "0000101101101000" =>
						DD(31, 36) <= packet_in;
						counter <= "0000101101101001";
						WHEN "0000101101101001" =>
						DD(31, 37) <= packet_in;
						counter <= "0000101101101010";
						WHEN "0000101101101010" =>
						DD(31, 38) <= packet_in;
						counter <= "0000101101101011";
						WHEN "0000101101101011" =>
						DD(31, 39) <= packet_in;
						counter <= "0000101101101100";
						WHEN "0000101101101100" =>
						DD(31, 40) <= packet_in;
						counter <= "0000101101101101";
						WHEN "0000101101101101" =>
						DD(31, 41) <= packet_in;
						counter <= "0000101101101110";
						WHEN "0000101101101110" =>
						DD(31, 42) <= packet_in;
						counter <= "0000101101101111";
						WHEN "0000101101101111" =>
						DD(31, 43) <= packet_in;
						counter <= "0000101101110000";
						WHEN "0000101101110000" =>
						DD(31, 44) <= packet_in;
						counter <= "0000101101110001";
						WHEN "0000101101110001" =>
						DD(31, 45) <= packet_in;
						counter <= "0000101101110010";
						WHEN "0000101101110010" =>
						DD(31, 46) <= packet_in;
						counter <= "0000101101110011";
						WHEN "0000101101110011" =>
						DD(31, 47) <= packet_in;
						counter <= "0000101101110100";
						WHEN "0000101101110100" =>
						DD(31, 48) <= packet_in;
						counter <= "0000101101110101";
						WHEN "0000101101110101" =>
						DD(31, 49) <= packet_in;
						counter <= "0000101101110110";
						WHEN "0000101101110110" =>
						DD(31, 50) <= packet_in;
						counter <= "0000101101110111";
						WHEN "0000101101110111" =>
						DD(31, 51) <= packet_in;
						counter <= "0000101101111000";
						WHEN "0000101101111000" =>
						DD(31, 52) <= packet_in;
						counter <= "0000101101111001";
						WHEN "0000101101111001" =>
						DD(31, 53) <= packet_in;
						counter <= "0000101101111010";
						WHEN "0000101101111010" =>
						DD(31, 54) <= packet_in;
						counter <= "0000101101111011";
						WHEN "0000101101111011" =>
						DD(31, 55) <= packet_in;
						counter <= "0000101101111100";
						WHEN "0000101101111100" =>
						DD(31, 56) <= packet_in;
						counter <= "0000101101111101";
						WHEN "0000101101111101" =>
						DD(31, 57) <= packet_in;
						counter <= "0000101101111110";
						WHEN "0000101101111110" =>
						DD(31, 58) <= packet_in;
						counter <= "0000101101111111";
						WHEN "0000101101111111" =>
						DD(31, 59) <= packet_in;
						counter <= "0000101110000000";
						WHEN "0000101110000000" =>
						DD(31, 60) <= packet_in;
						counter <= "0000101110000001";
						WHEN "0000101110000001" =>
						DD(31, 61) <= packet_in;
						counter <= "0000101110000010";
						WHEN "0000101110000010" =>
						DD(31, 62) <= packet_in;
						counter <= "0000101110000011";
						WHEN "0000101110000011" =>
						DD(31, 63) <= packet_in;
						counter <= "0000101110000100";
						WHEN "0000101110000100" =>
						DD(31, 64) <= packet_in;
						counter <= "0000101110000101";
						WHEN "0000101110000101" =>
						DD(31, 65) <= packet_in;
						counter <= "0000101110000110";
						WHEN "0000101110000110" =>
						DD(31, 66) <= packet_in;
						counter <= "0000101110000111";
						WHEN "0000101110000111" =>
						DD(31, 67) <= packet_in;
						counter <= "0000101110001000";
						WHEN "0000101110001000" =>
						DD(31, 68) <= packet_in;
						counter <= "0000101110001001";
						WHEN "0000101110001001" =>
						DD(31, 69) <= packet_in;
						counter <= "0000101110001010";
						WHEN "0000101110001010" =>
						DD(31, 70) <= packet_in;
						counter <= "0000101110001011";
						WHEN "0000101110001011" =>
						DD(31, 71) <= packet_in;
						counter <= "0000101110001100";
						WHEN "0000101110001100" =>
						DD(31, 72) <= packet_in;
						counter <= "0000101110001101";
						WHEN "0000101110001101" =>
						DD(31, 73) <= packet_in;
						counter <= "0000101110001110";
						WHEN "0000101110001110" =>
						DD(31, 74) <= packet_in;
						counter <= "0000101110001111";
						WHEN "0000101110001111" =>
						DD(31, 75) <= packet_in;
						counter <= "0000101110010000";
						WHEN "0000101110010000" =>
						DD(31, 76) <= packet_in;
						counter <= "0000101110010001";
						WHEN "0000101110010001" =>
						DD(31, 77) <= packet_in;
						counter <= "0000101110010010";
						WHEN "0000101110010010" =>
						DD(31, 78) <= packet_in;
						counter <= "0000101110010011";
						WHEN "0000101110010011" =>
						DD(31, 79) <= packet_in;
						counter <= "0000101110010100";
						WHEN "0000101110010100" =>
						DD(31, 80) <= packet_in;
						counter <= "0000101110010101";
						WHEN "0000101110010101" =>
						DD(31, 81) <= packet_in;
						counter <= "0000101110010110";
						WHEN "0000101110010110" =>
						DD(31, 82) <= packet_in;
						counter <= "0000101110010111";
						WHEN "0000101110010111" =>
						DD(31, 83) <= packet_in;
						counter <= "0000101110011000";
						WHEN "0000101110011000" =>
						DD(31, 84) <= packet_in;
						counter <= "0000101110011001";
						WHEN "0000101110011001" =>
						DD(31, 85) <= packet_in;
						counter <= "0000101110011010";
						WHEN "0000101110011010" =>
						DD(31, 86) <= packet_in;
						counter <= "0000101110011011";
						WHEN "0000101110011011" =>
						DD(31, 87) <= packet_in;
						counter <= "0000101110011100";
						WHEN "0000101110011100" =>
						DD(31, 88) <= packet_in;
						counter <= "0000101110011101";
						WHEN "0000101110011101" =>
						DD(31, 89) <= packet_in;
						counter <= "0000101110011110";
						WHEN "0000101110011110" =>
						DD(31, 90) <= packet_in;
						counter <= "0000101110011111";
						WHEN "0000101110011111" =>
						DD(31, 91) <= packet_in;
						counter <= "0000000000000000";
						dd_received <= '1';
--						WHEN "0000101110100000" =>
						
						WHEN OTHERS =>
						NULL;
					END CASE;

					WHEN OTHERS =>
					NULL;
				END CASE;
			else
				dd_received <= '0';
				hello_received <= '0';
			END IF;
		END IF;
	END PROCESS;

--process(hello_done)
--begin
--	hello_received <= '1';
--end process;

END packetParser_arc;