-- TestBench Template 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.main_package.ALL;

ENTITY testbench IS
END testbench;

ARCHITECTURE behavior OF testbench IS

	COMPONENT main_OSPF IS
		PORT (
			-- input packets
			-- valid_i will be 1 if packet_i is coming
			packet_in1 : IN std_logic_vector(7 DOWNTO 0);
			packet_in2 : IN std_logic_vector(7 DOWNTO 0);
			packet_in3 : IN std_logic_vector(7 DOWNTO 0);
			packet_in4 : IN std_logic_vector(7 DOWNTO 0);
			packet_in5 : IN std_logic_vector(7 DOWNTO 0);
			packet_in6 : IN std_logic_vector(7 DOWNTO 0);
			packet_in7 : IN std_logic_vector(7 DOWNTO 0);
			packet_in8 : IN std_logic_vector(7 DOWNTO 0);
			valid_in1 : IN std_logic;
			valid_in2 : IN std_logic;
			valid_in3 : IN std_logic;
			valid_in4 : IN std_logic;
			valid_in5 : IN std_logic;
			valid_in6 : IN std_logic;
			valid_in7 : IN std_logic;
			valid_in8 : IN std_logic;

			-- clocks to be decided according to needs
			clk : IN std_logic;
			-- clocks end here
			-- output packets
			gateway_ip : OUT ip_addr_array;
			gateway_node : OUT RAM_FOR_NEXTHOP;
			packet_out1 : OUT std_logic_vector(7 DOWNTO 0);
			packet_out2 : OUT std_logic_vector(7 DOWNTO 0);
			packet_out3 : OUT std_logic_vector(7 DOWNTO 0);
			packet_out4 : OUT std_logic_vector(7 DOWNTO 0);
			packet_out5 : OUT std_logic_vector(7 DOWNTO 0);
			packet_out6 : OUT std_logic_vector(7 DOWNTO 0);
			packet_out7 : OUT std_logic_vector(7 DOWNTO 0);
			packet_out8 : OUT std_logic_vector(7 DOWNTO 0);
			valid_out1 : OUT std_logic;
			valid_out2 : OUT std_logic;
			valid_out3 : OUT std_logic;
			valid_out4 : OUT std_logic;
			valid_out5 : OUT std_logic;
			valid_out6 : OUT std_logic;
			valid_out7 : OUT std_logic;
			valid_out8 : OUT std_logic);
	END COMPONENT main_OSPF;

	SIGNAL packet_in1 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL packet_in2 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL packet_in3 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL packet_in4 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL packet_in5 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL packet_in6 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL packet_in7 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL packet_in8 : std_logic_vector(7 DOWNTO 0) := "00000000";
	SIGNAL valid_in1 : std_logic := '0';
	SIGNAL valid_in2 : std_logic := '0';
	SIGNAL valid_in3 : std_logic := '0';
	SIGNAL valid_in4 : std_logic := '0';
	SIGNAL valid_in5 : std_logic := '0';
	SIGNAL valid_in6 : std_logic := '0';
	SIGNAL valid_in7 : std_logic := '0';
	SIGNAL valid_in8 : std_logic := '0';

	-- clocks to be decided according to needs
	SIGNAL clk : std_logic := '0';
	SIGNAL gateway_ip : ip_addr_array;
	SIGNAL gateway_node : RAM_FOR_NEXTHOP;
	SIGNAL packet_out1 : std_logic_vector(7 DOWNTO 0);
	SIGNAL packet_out2 : std_logic_vector(7 DOWNTO 0);
	SIGNAL packet_out3 : std_logic_vector(7 DOWNTO 0);
	SIGNAL packet_out4 : std_logic_vector(7 DOWNTO 0);
	SIGNAL packet_out5 : std_logic_vector(7 DOWNTO 0);
	SIGNAL packet_out6 : std_logic_vector(7 DOWNTO 0);
	SIGNAL packet_out7 : std_logic_vector(7 DOWNTO 0);
	SIGNAL packet_out8 : std_logic_vector(7 DOWNTO 0);
	SIGNAL valid_out1 : std_logic;
	SIGNAL valid_out2 : std_logic;
	SIGNAL valid_out3 : std_logic;
	SIGNAL valid_out4 : std_logic;
	SIGNAL valid_out5 : std_logic;
	SIGNAL valid_out6 : std_logic;
	SIGNAL valid_out7 : std_logic;
	SIGNAL valid_out8 : std_logic;

	CONSTANT clk_period : TIME := 1 ns;
BEGIN

	-- Component Instantiation
	uut : main_OSPF PORT MAP(
		-- valid_i will be 1 if packet_i is coming
		packet_in1,
		packet_in2,
		packet_in3,
		packet_in4,
		packet_in5,
		packet_in6,
		packet_in7,
		packet_in8,
		valid_in1,
		valid_in2,
		valid_in3,
		valid_in4,
		valid_in5,
		valid_in6,
		valid_in7,
		valid_in8,
		clk,
		gateway_ip,
		gateway_node,
		packet_out1,
		packet_out2,
		packet_out3,
		packet_out4,
		packet_out5,
		packet_out6,
		packet_out7,
		packet_out8,
		valid_out1,
		valid_out2,
		valid_out3,
		valid_out4,
		valid_out5,
		valid_out6,
		valid_out7,
		valid_out8);

	clk_process : PROCESS
	BEGIN
		clk <= '0';
		WAIT FOR clk_period/2;
		clk <= '1';
		WAIT FOR clk_period/2;
	END PROCESS;
	--  Test Bench Statements
	tb : PROCESS
	BEGIN
		WAIT FOR 10 ns;
		valid_in1 <= '1';
		valid_in2 <= '1';
		valid_in3 <= '1';
		valid_in4 <= '1';
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		-- I/P for PACKET TYPE
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		-- I/P for PACKET LENGTH
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for ROUTER ID
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for AREA ID
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for CHECKSUM
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for AU TYPE
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for AUTHENTICATION
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for NETWORK MASK
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for HELLO INTERVAL
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for OPTIONS
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for RTE PRI
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for ROUTER DEAD INTERVAL
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Designated ROUTER
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for BACKUP ROUTER
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour0
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour1
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in4 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in1 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour2
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour3
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour4
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour5
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour6
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		-- I/P for Neighbour7
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		--  wait for clk_period;
		--  wait for clk_period;
		valid_in1 <= '0'; 
		valid_in2 <= '0'; 
		valid_in3 <= '0';
		valid_in4 <= '0'; 
		WAIT FOR 20 ns;
		valid_in1 <= '1';
		valid_in2 <= '1';
		valid_in3 <= '1';
		valid_in4 <= '1';
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00001011";
		packet_in2 <= "00001011";
		packet_in3 <= "00001011";
		packet_in4 <= "00001011";
		WAIT FOR clk_period;
		packet_in1 <= "10001100";
		packet_in2 <= "10001100";
		packet_in3 <= "10001100";
		packet_in4 <= "10001100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001100";
		packet_in2 <= "00001100";
		packet_in3 <= "00001100";
		packet_in4 <= "00001100";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001100";
		packet_in2 <= "00001100";
		packet_in3 <= "00001100";
		packet_in4 <= "00001100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001001";
		packet_in2 <= "00001001";
		packet_in3 <= "00001001";
		packet_in4 <= "00001001";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001001";
		packet_in2 <= "00001001";
		packet_in3 <= "00001001";
		packet_in4 <= "00001001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000111";
		packet_in2 <= "00000111";
		packet_in3 <= "00000111";
		packet_in4 <= "00000111";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000111";
		packet_in2 <= "00000111";
		packet_in3 <= "00000111";
		packet_in4 <= "00000111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000111";
		packet_in2 <= "00000111";
		packet_in3 <= "00000111";
		packet_in4 <= "00000111";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000111";
		packet_in2 <= "00000111";
		packet_in3 <= "00000111";
		packet_in4 <= "00000111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000111";
		packet_in2 <= "00000111";
		packet_in3 <= "00000111";
		packet_in4 <= "00000111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000111";
		packet_in2 <= "00000111";
		packet_in3 <= "00000111";
		packet_in4 <= "00000111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000100";
		packet_in2 <= "00000100";
		packet_in3 <= "00000100";
		packet_in4 <= "00000100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001000";
		packet_in2 <= "00001000";
		packet_in3 <= "00001000";
		packet_in4 <= "00001000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001000";
		packet_in2 <= "00001000";
		packet_in3 <= "00001000";
		packet_in4 <= "00001000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001010";
		packet_in2 <= "00001010";
		packet_in3 <= "00001010";
		packet_in4 <= "00001010";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001010";
		packet_in2 <= "00001010";
		packet_in3 <= "00001010";
		packet_in4 <= "00001010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001011";
		packet_in2 <= "00001011";
		packet_in3 <= "00001011";
		packet_in4 <= "00001011";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001011";
		packet_in2 <= "00001011";
		packet_in3 <= "00001011";
		packet_in4 <= "00001011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001001";
		packet_in2 <= "00001001";
		packet_in3 <= "00001001";
		packet_in4 <= "00001001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001001";
		packet_in2 <= "00001001";
		packet_in3 <= "00001001";
		packet_in4 <= "00001001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001100";
		packet_in2 <= "00001100";
		packet_in3 <= "00001100";
		packet_in4 <= "00001100";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001100";
		packet_in2 <= "00001100";
		packet_in3 <= "00001100";
		packet_in4 <= "00001100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001010";
		packet_in2 <= "00001010";
		packet_in3 <= "00001010";
		packet_in4 <= "00001010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001010";
		packet_in2 <= "00001010";
		packet_in3 <= "00001010";
		packet_in4 <= "00001010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001000";
		packet_in2 <= "00001000";
		packet_in3 <= "00001000";
		packet_in4 <= "00001000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001000";
		packet_in2 <= "00001000";
		packet_in3 <= "00001000";
		packet_in4 <= "00001000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000110";
		packet_in2 <= "00000110";
		packet_in3 <= "00000110";
		packet_in4 <= "00000110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001011";
		packet_in2 <= "00001011";
		packet_in3 <= "00001011";
		packet_in4 <= "00001011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001011";
		packet_in2 <= "00001011";
		packet_in3 <= "00001011";
		packet_in4 <= "00001011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001000";
		packet_in2 <= "00001000";
		packet_in3 <= "00001000";
		packet_in4 <= "00001000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001000";
		packet_in2 <= "00001000";
		packet_in3 <= "00001000";
		packet_in4 <= "00001000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001100";
		packet_in2 <= "00001100";
		packet_in3 <= "00001100";
		packet_in4 <= "00001100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001100";
		packet_in2 <= "00001100";
		packet_in3 <= "00001100";
		packet_in4 <= "00001100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001001";
		packet_in2 <= "00001001";
		packet_in3 <= "00001001";
		packet_in4 <= "00001001";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001001";
		packet_in2 <= "00001001";
		packet_in3 <= "00001001";
		packet_in4 <= "00001001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001101";
		packet_in2 <= "00001101";
		packet_in3 <= "00001101";
		packet_in4 <= "00001101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001010";
		packet_in2 <= "00001010";
		packet_in3 <= "00001010";
		packet_in4 <= "00001010";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001010";
		packet_in2 <= "00001010";
		packet_in3 <= "00001010";
		packet_in4 <= "00001010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001011";
		packet_in2 <= "00001011";
		packet_in3 <= "00001011";
		packet_in4 <= "00001011";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001011";
		packet_in2 <= "00001011";
		packet_in3 <= "00001011";
		packet_in4 <= "00001011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001110";
		packet_in2 <= "00001110";
		packet_in3 <= "00001110";
		packet_in4 <= "00001110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000101";
		packet_in2 <= "00000101";
		packet_in3 <= "00000101";
		packet_in4 <= "00000101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000011";
		packet_in2 <= "00000011";
		packet_in3 <= "00000011";
		packet_in4 <= "00000011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000010";
		packet_in2 <= "00000010";
		packet_in3 <= "00000010";
		packet_in4 <= "00000010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00001111";
		packet_in2 <= "00001111";
		packet_in3 <= "00001111";
		packet_in4 <= "00001111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00001111";
		packet_in2 <= "00001111";
		packet_in3 <= "00001111";
		packet_in4 <= "00001111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010000";
		packet_in2 <= "00010000";
		packet_in3 <= "00010000";
		packet_in4 <= "00010000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010000";
		packet_in2 <= "00010000";
		packet_in3 <= "00010000";
		packet_in4 <= "00010000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010001";
		packet_in2 <= "00010001";
		packet_in3 <= "00010001";
		packet_in4 <= "00010001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010001";
		packet_in2 <= "00010001";
		packet_in3 <= "00010001";
		packet_in4 <= "00010001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010010";
		packet_in2 <= "00010010";
		packet_in3 <= "00010010";
		packet_in4 <= "00010010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010010";
		packet_in2 <= "00010010";
		packet_in3 <= "00010010";
		packet_in4 <= "00010010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010011";
		packet_in2 <= "00010011";
		packet_in3 <= "00010011";
		packet_in4 <= "00010011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010011";
		packet_in2 <= "00010011";
		packet_in3 <= "00010011";
		packet_in4 <= "00010011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010100";
		packet_in2 <= "00010100";
		packet_in3 <= "00010100";
		packet_in4 <= "00010100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010100";
		packet_in2 <= "00010100";
		packet_in3 <= "00010100";
		packet_in4 <= "00010100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010101";
		packet_in2 <= "00010101";
		packet_in3 <= "00010101";
		packet_in4 <= "00010101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010101";
		packet_in2 <= "00010101";
		packet_in3 <= "00010101";
		packet_in4 <= "00010101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010110";
		packet_in2 <= "00010110";
		packet_in3 <= "00010110";
		packet_in4 <= "00010110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010110";
		packet_in2 <= "00010110";
		packet_in3 <= "00010110";
		packet_in4 <= "00010110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00010111";
		packet_in2 <= "00010111";
		packet_in3 <= "00010111";
		packet_in4 <= "00010111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00010111";
		packet_in2 <= "00010111";
		packet_in3 <= "00010111";
		packet_in4 <= "00010111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011000";
		packet_in2 <= "00011000";
		packet_in3 <= "00011000";
		packet_in4 <= "00011000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011000";
		packet_in2 <= "00011000";
		packet_in3 <= "00011000";
		packet_in4 <= "00011000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011001";
		packet_in2 <= "00011001";
		packet_in3 <= "00011001";
		packet_in4 <= "00011001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011001";
		packet_in2 <= "00011001";
		packet_in3 <= "00011001";
		packet_in4 <= "00011001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011010";
		packet_in2 <= "00011010";
		packet_in3 <= "00011010";
		packet_in4 <= "00011010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011010";
		packet_in2 <= "00011010";
		packet_in3 <= "00011010";
		packet_in4 <= "00011010";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011011";
		packet_in2 <= "00011011";
		packet_in3 <= "00011011";
		packet_in4 <= "00011011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011011";
		packet_in2 <= "00011011";
		packet_in3 <= "00011011";
		packet_in4 <= "00011011";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011100";
		packet_in2 <= "00011100";
		packet_in3 <= "00011100";
		packet_in4 <= "00011100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011100";
		packet_in2 <= "00011100";
		packet_in3 <= "00011100";
		packet_in4 <= "00011100";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011101";
		packet_in2 <= "00011101";
		packet_in3 <= "00011101";
		packet_in4 <= "00011101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011101";
		packet_in2 <= "00011101";
		packet_in3 <= "00011101";
		packet_in4 <= "00011101";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011110";
		packet_in2 <= "00011110";
		packet_in3 <= "00011110";
		packet_in4 <= "00011110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011110";
		packet_in2 <= "00011110";
		packet_in3 <= "00011110";
		packet_in4 <= "00011110";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00011111";
		packet_in2 <= "00011111";
		packet_in3 <= "00011111";
		packet_in4 <= "00011111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00011111";
		packet_in2 <= "00011111";
		packet_in3 <= "00011111";
		packet_in4 <= "00011111";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000001";
		packet_in2 <= "00000001";
		packet_in3 <= "00000001";
		packet_in4 <= "00000001";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "11000000";
		packet_in2 <= "11000000";
		packet_in3 <= "11000000";
		packet_in4 <= "11000000";
		WAIT FOR clk_period;
		packet_in1 <= "10101000";
		packet_in2 <= "10101000";
		packet_in3 <= "10101000";
		packet_in4 <= "10101000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		packet_in1 <= "00000000";
		packet_in2 <= "00000000";
		packet_in3 <= "00000000";
		packet_in4 <= "00000000";
		WAIT FOR clk_period;
		valid_in1 <= '0';
		valid_in2 <= '0';
		valid_in3 <= '0';
		valid_in4 <= '0';
		WAIT FOR 20 ns;
		WAIT; -- will wait forever
	END PROCESS tb;
	--  End Test Bench 

END;