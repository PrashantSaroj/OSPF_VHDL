LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.numeric_std.ALL;
USE WORK.main_package.ALL;

ENTITY extract_info IS
	PORT (
		control : in std_logic;
		DD : IN databaseDescription;
		graph : OUT RAM_FOR_GRAPH;
		IP_ADDR : OUT ip_addr_array;
		extraction_done: out std_logic);
END extract_info;

ARCHITECTURE behavioural OF extract_info IS

BEGIN
	-- assumption router ids are 0-31
	process(control) is 

	VARIABLE d1, d2, d3, d4 : std_logic_vector(7 DOWNTO 0):="00000000";
	VARIABLE e1, e2, e3, e4 : std_logic_vector(7 DOWNTO 0):="00000000";
	VARIABLE d, e : std_logic_vector(31 DOWNTO 0):="00000000000000000000000000000000";

	begin
	if control = '1' then 
	d1 := DD(0, 4);
			d2 := DD(0, 5);
			d3 := DD(0, 6);
			d4 := DD(0, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(0, 0);
			e2 := DD(0, 1);
			e3 := DD(0, 2);
			e4 := DD(0, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(1, 4);
			d2 := DD(1, 5);
			d3 := DD(1, 6);
			d4 := DD(1, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(1, 0);
			e2 := DD(1, 1);
			e3 := DD(1, 2);
			e4 := DD(1, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(2, 4);
			d2 := DD(2, 5);
			d3 := DD(2, 6);
			d4 := DD(2, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(2, 0);
			e2 := DD(2, 1);
			e3 := DD(2, 2);
			e4 := DD(2, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(3, 4);
			d2 := DD(3, 5);
			d3 := DD(3, 6);
			d4 := DD(3, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(3, 0);
			e2 := DD(3, 1);
			e3 := DD(3, 2);
			e4 := DD(3, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(4, 4);
			d2 := DD(4, 5);
			d3 := DD(4, 6);
			d4 := DD(4, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(4, 0);
			e2 := DD(4, 1);
			e3 := DD(4, 2);
			e4 := DD(4, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(5, 4);
			d2 := DD(5, 5);
			d3 := DD(5, 6);
			d4 := DD(5, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(5, 0);
			e2 := DD(5, 1);
			e3 := DD(5, 2);
			e4 := DD(5, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(6, 4);
			d2 := DD(6, 5);
			d3 := DD(6, 6);
			d4 := DD(6, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(6, 0);
			e2 := DD(6, 1);
			e3 := DD(6, 2);
			e4 := DD(6, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(7, 4);
			d2 := DD(7, 5);
			d3 := DD(7, 6);
			d4 := DD(7, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(7, 0);
			e2 := DD(7, 1);
			e3 := DD(7, 2);
			e4 := DD(7, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(8, 4);
			d2 := DD(8, 5);
			d3 := DD(8, 6);
			d4 := DD(8, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(8, 0);
			e2 := DD(8, 1);
			e3 := DD(8, 2);
			e4 := DD(8, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(9, 4);
			d2 := DD(9, 5);
			d3 := DD(9, 6);
			d4 := DD(9, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(9, 0);
			e2 := DD(9, 1);
			e3 := DD(9, 2);
			e4 := DD(9, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(10, 4);
			d2 := DD(10, 5);
			d3 := DD(10, 6);
			d4 := DD(10, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(10, 0);
			e2 := DD(10, 1);
			e3 := DD(10, 2);
			e4 := DD(10, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(11, 4);
			d2 := DD(11, 5);
			d3 := DD(11, 6);
			d4 := DD(11, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(11, 0);
			e2 := DD(11, 1);
			e3 := DD(11, 2);
			e4 := DD(11, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(12, 4);
			d2 := DD(12, 5);
			d3 := DD(12, 6);
			d4 := DD(12, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(12, 0);
			e2 := DD(12, 1);
			e3 := DD(12, 2);
			e4 := DD(12, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(13, 4);
			d2 := DD(13, 5);
			d3 := DD(13, 6);
			d4 := DD(13, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(13, 0);
			e2 := DD(13, 1);
			e3 := DD(13, 2);
			e4 := DD(13, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(14, 4);
			d2 := DD(14, 5);
			d3 := DD(14, 6);
			d4 := DD(14, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(14, 0);
			e2 := DD(14, 1);
			e3 := DD(14, 2);
			e4 := DD(14, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(15, 4);
			d2 := DD(15, 5);
			d3 := DD(15, 6);
			d4 := DD(15, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(15, 0);
			e2 := DD(15, 1);
			e3 := DD(15, 2);
			e4 := DD(15, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(16, 4);
			d2 := DD(16, 5);
			d3 := DD(16, 6);
			d4 := DD(16, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(16, 0);
			e2 := DD(16, 1);
			e3 := DD(16, 2);
			e4 := DD(16, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(17, 4);
			d2 := DD(17, 5);
			d3 := DD(17, 6);
			d4 := DD(17, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(17, 0);
			e2 := DD(17, 1);
			e3 := DD(17, 2);
			e4 := DD(17, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(18, 4);
			d2 := DD(18, 5);
			d3 := DD(18, 6);
			d4 := DD(18, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(18, 0);
			e2 := DD(18, 1);
			e3 := DD(18, 2);
			e4 := DD(18, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(19, 4);
			d2 := DD(19, 5);
			d3 := DD(19, 6);
			d4 := DD(19, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(19, 0);
			e2 := DD(19, 1);
			e3 := DD(19, 2);
			e4 := DD(19, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(20, 4);
			d2 := DD(20, 5);
			d3 := DD(20, 6);
			d4 := DD(20, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(20, 0);
			e2 := DD(20, 1);
			e3 := DD(20, 2);
			e4 := DD(20, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(21, 4);
			d2 := DD(21, 5);
			d3 := DD(21, 6);
			d4 := DD(21, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(21, 0);
			e2 := DD(21, 1);
			e3 := DD(21, 2);
			e4 := DD(21, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(22, 4);
			d2 := DD(22, 5);
			d3 := DD(22, 6);
			d4 := DD(22, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(22, 0);
			e2 := DD(22, 1);
			e3 := DD(22, 2);
			e4 := DD(22, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(23, 4);
			d2 := DD(23, 5);
			d3 := DD(23, 6);
			d4 := DD(23, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(23, 0);
			e2 := DD(23, 1);
			e3 := DD(23, 2);
			e4 := DD(23, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(24, 4);
			d2 := DD(24, 5);
			d3 := DD(24, 6);
			d4 := DD(24, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(24, 0);
			e2 := DD(24, 1);
			e3 := DD(24, 2);
			e4 := DD(24, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(25, 4);
			d2 := DD(25, 5);
			d3 := DD(25, 6);
			d4 := DD(25, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(25, 0);
			e2 := DD(25, 1);
			e3 := DD(25, 2);
			e4 := DD(25, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(26, 4);
			d2 := DD(26, 5);
			d3 := DD(26, 6);
			d4 := DD(26, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(26, 0);
			e2 := DD(26, 1);
			e3 := DD(26, 2);
			e4 := DD(26, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(27, 4);
			d2 := DD(27, 5);
			d3 := DD(27, 6);
			d4 := DD(27, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(27, 0);
			e2 := DD(27, 1);
			e3 := DD(27, 2);
			e4 := DD(27, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(28, 4);
			d2 := DD(28, 5);
			d3 := DD(28, 6);
			d4 := DD(28, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(28, 0);
			e2 := DD(28, 1);
			e3 := DD(28, 2);
			e4 := DD(28, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(29, 4);
			d2 := DD(29, 5);
			d3 := DD(29, 6);
			d4 := DD(29, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(29, 0);
			e2 := DD(29, 1);
			e3 := DD(29, 2);
			e4 := DD(29, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(30, 4);
			d2 := DD(30, 5);
			d3 := DD(30, 6);
			d4 := DD(30, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(30, 0);
			e2 := DD(30, 1);
			e3 := DD(30, 2);
			e4 := DD(30, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
			d1 := DD(31, 4);
			d2 := DD(31, 5);
			d3 := DD(31, 6);
			d4 := DD(31, 7);
			d := d1 & d2 & d3 & d4;
			e1 := DD(31, 0);
			e2 := DD(31, 1);
			e3 := DD(31, 2);
			e4 := DD(31, 3);
			e := e1 & e2 & e3 & e4;
			IP_ADDR(to_integer(unsigned(d))) <= e;
		-- initialize cost to maximum
		graph(0,0) <= "11111111";
		graph(0,1) <= "11111111";
		graph(0,2) <= "11111111";
		graph(0,3) <= "11111111";
		graph(0,4) <= "11111111";
		graph(0,5) <= "11111111";
		graph(0,6) <= "11111111";
		graph(0,7) <= "11111111";
		graph(0,8) <= "11111111";
		graph(0,9) <= "11111111";
		graph(0,10) <= "11111111";
		graph(0,11) <= "11111111";
		graph(0,12) <= "11111111";
		graph(0,13) <= "11111111";
		graph(0,14) <= "11111111";
		graph(0,15) <= "11111111";
		graph(0,16) <= "11111111";
		graph(0,17) <= "11111111";
		graph(0,18) <= "11111111";
		graph(0,19) <= "11111111";
		graph(0,20) <= "11111111";
		graph(0,21) <= "11111111";
		graph(0,22) <= "11111111";
		graph(0,23) <= "11111111";
		graph(0,24) <= "11111111";
		graph(0,25) <= "11111111";
		graph(0,26) <= "11111111";
		graph(0,27) <= "11111111";
		graph(0,28) <= "11111111";
		graph(0,29) <= "11111111";
		graph(0,30) <= "11111111";
		graph(0,31) <= "11111111";
		graph(1,0) <= "11111111";
		graph(1,1) <= "11111111";
		graph(1,2) <= "11111111";
		graph(1,3) <= "11111111";
		graph(1,4) <= "11111111";
		graph(1,5) <= "11111111";
		graph(1,6) <= "11111111";
		graph(1,7) <= "11111111";
		graph(1,8) <= "11111111";
		graph(1,9) <= "11111111";
		graph(1,10) <= "11111111";
		graph(1,11) <= "11111111";
		graph(1,12) <= "11111111";
		graph(1,13) <= "11111111";
		graph(1,14) <= "11111111";
		graph(1,15) <= "11111111";
		graph(1,16) <= "11111111";
		graph(1,17) <= "11111111";
		graph(1,18) <= "11111111";
		graph(1,19) <= "11111111";
		graph(1,20) <= "11111111";
		graph(1,21) <= "11111111";
		graph(1,22) <= "11111111";
		graph(1,23) <= "11111111";
		graph(1,24) <= "11111111";
		graph(1,25) <= "11111111";
		graph(1,26) <= "11111111";
		graph(1,27) <= "11111111";
		graph(1,28) <= "11111111";
		graph(1,29) <= "11111111";
		graph(1,30) <= "11111111";
		graph(1,31) <= "11111111";
		graph(2,0) <= "11111111";
		graph(2,1) <= "11111111";
		graph(2,2) <= "11111111";
		graph(2,3) <= "11111111";
		graph(2,4) <= "11111111";
		graph(2,5) <= "11111111";
		graph(2,6) <= "11111111";
		graph(2,7) <= "11111111";
		graph(2,8) <= "11111111";
		graph(2,9) <= "11111111";
		graph(2,10) <= "11111111";
		graph(2,11) <= "11111111";
		graph(2,12) <= "11111111";
		graph(2,13) <= "11111111";
		graph(2,14) <= "11111111";
		graph(2,15) <= "11111111";
		graph(2,16) <= "11111111";
		graph(2,17) <= "11111111";
		graph(2,18) <= "11111111";
		graph(2,19) <= "11111111";
		graph(2,20) <= "11111111";
		graph(2,21) <= "11111111";
		graph(2,22) <= "11111111";
		graph(2,23) <= "11111111";
		graph(2,24) <= "11111111";
		graph(2,25) <= "11111111";
		graph(2,26) <= "11111111";
		graph(2,27) <= "11111111";
		graph(2,28) <= "11111111";
		graph(2,29) <= "11111111";
		graph(2,30) <= "11111111";
		graph(2,31) <= "11111111";
		graph(3,0) <= "11111111";
		graph(3,1) <= "11111111";
		graph(3,2) <= "11111111";
		graph(3,3) <= "11111111";
		graph(3,4) <= "11111111";
		graph(3,5) <= "11111111";
		graph(3,6) <= "11111111";
		graph(3,7) <= "11111111";
		graph(3,8) <= "11111111";
		graph(3,9) <= "11111111";
		graph(3,10) <= "11111111";
		graph(3,11) <= "11111111";
		graph(3,12) <= "11111111";
		graph(3,13) <= "11111111";
		graph(3,14) <= "11111111";
		graph(3,15) <= "11111111";
		graph(3,16) <= "11111111";
		graph(3,17) <= "11111111";
		graph(3,18) <= "11111111";
		graph(3,19) <= "11111111";
		graph(3,20) <= "11111111";
		graph(3,21) <= "11111111";
		graph(3,22) <= "11111111";
		graph(3,23) <= "11111111";
		graph(3,24) <= "11111111";
		graph(3,25) <= "11111111";
		graph(3,26) <= "11111111";
		graph(3,27) <= "11111111";
		graph(3,28) <= "11111111";
		graph(3,29) <= "11111111";
		graph(3,30) <= "11111111";
		graph(3,31) <= "11111111";
		graph(4,0) <= "11111111";
		graph(4,1) <= "11111111";
		graph(4,2) <= "11111111";
		graph(4,3) <= "11111111";
		graph(4,4) <= "11111111";
		graph(4,5) <= "11111111";
		graph(4,6) <= "11111111";
		graph(4,7) <= "11111111";
		graph(4,8) <= "11111111";
		graph(4,9) <= "11111111";
		graph(4,10) <= "11111111";
		graph(4,11) <= "11111111";
		graph(4,12) <= "11111111";
		graph(4,13) <= "11111111";
		graph(4,14) <= "11111111";
		graph(4,15) <= "11111111";
		graph(4,16) <= "11111111";
		graph(4,17) <= "11111111";
		graph(4,18) <= "11111111";
		graph(4,19) <= "11111111";
		graph(4,20) <= "11111111";
		graph(4,21) <= "11111111";
		graph(4,22) <= "11111111";
		graph(4,23) <= "11111111";
		graph(4,24) <= "11111111";
		graph(4,25) <= "11111111";
		graph(4,26) <= "11111111";
		graph(4,27) <= "11111111";
		graph(4,28) <= "11111111";
		graph(4,29) <= "11111111";
		graph(4,30) <= "11111111";
		graph(4,31) <= "11111111";
		graph(5,0) <= "11111111";
		graph(5,1) <= "11111111";
		graph(5,2) <= "11111111";
		graph(5,3) <= "11111111";
		graph(5,4) <= "11111111";
		graph(5,5) <= "11111111";
		graph(5,6) <= "11111111";
		graph(5,7) <= "11111111";
		graph(5,8) <= "11111111";
		graph(5,9) <= "11111111";
		graph(5,10) <= "11111111";
		graph(5,11) <= "11111111";
		graph(5,12) <= "11111111";
		graph(5,13) <= "11111111";
		graph(5,14) <= "11111111";
		graph(5,15) <= "11111111";
		graph(5,16) <= "11111111";
		graph(5,17) <= "11111111";
		graph(5,18) <= "11111111";
		graph(5,19) <= "11111111";
		graph(5,20) <= "11111111";
		graph(5,21) <= "11111111";
		graph(5,22) <= "11111111";
		graph(5,23) <= "11111111";
		graph(5,24) <= "11111111";
		graph(5,25) <= "11111111";
		graph(5,26) <= "11111111";
		graph(5,27) <= "11111111";
		graph(5,28) <= "11111111";
		graph(5,29) <= "11111111";
		graph(5,30) <= "11111111";
		graph(5,31) <= "11111111";
		graph(6,0) <= "11111111";
		graph(6,1) <= "11111111";
		graph(6,2) <= "11111111";
		graph(6,3) <= "11111111";
		graph(6,4) <= "11111111";
		graph(6,5) <= "11111111";
		graph(6,6) <= "11111111";
		graph(6,7) <= "11111111";
		graph(6,8) <= "11111111";
		graph(6,9) <= "11111111";
		graph(6,10) <= "11111111";
		graph(6,11) <= "11111111";
		graph(6,12) <= "11111111";
		graph(6,13) <= "11111111";
		graph(6,14) <= "11111111";
		graph(6,15) <= "11111111";
		graph(6,16) <= "11111111";
		graph(6,17) <= "11111111";
		graph(6,18) <= "11111111";
		graph(6,19) <= "11111111";
		graph(6,20) <= "11111111";
		graph(6,21) <= "11111111";
		graph(6,22) <= "11111111";
		graph(6,23) <= "11111111";
		graph(6,24) <= "11111111";
		graph(6,25) <= "11111111";
		graph(6,26) <= "11111111";
		graph(6,27) <= "11111111";
		graph(6,28) <= "11111111";
		graph(6,29) <= "11111111";
		graph(6,30) <= "11111111";
		graph(6,31) <= "11111111";
		graph(7,0) <= "11111111";
		graph(7,1) <= "11111111";
		graph(7,2) <= "11111111";
		graph(7,3) <= "11111111";
		graph(7,4) <= "11111111";
		graph(7,5) <= "11111111";
		graph(7,6) <= "11111111";
		graph(7,7) <= "11111111";
		graph(7,8) <= "11111111";
		graph(7,9) <= "11111111";
		graph(7,10) <= "11111111";
		graph(7,11) <= "11111111";
		graph(7,12) <= "11111111";
		graph(7,13) <= "11111111";
		graph(7,14) <= "11111111";
		graph(7,15) <= "11111111";
		graph(7,16) <= "11111111";
		graph(7,17) <= "11111111";
		graph(7,18) <= "11111111";
		graph(7,19) <= "11111111";
		graph(7,20) <= "11111111";
		graph(7,21) <= "11111111";
		graph(7,22) <= "11111111";
		graph(7,23) <= "11111111";
		graph(7,24) <= "11111111";
		graph(7,25) <= "11111111";
		graph(7,26) <= "11111111";
		graph(7,27) <= "11111111";
		graph(7,28) <= "11111111";
		graph(7,29) <= "11111111";
		graph(7,30) <= "11111111";
		graph(7,31) <= "11111111";
		graph(8,0) <= "11111111";
		graph(8,1) <= "11111111";
		graph(8,2) <= "11111111";
		graph(8,3) <= "11111111";
		graph(8,4) <= "11111111";
		graph(8,5) <= "11111111";
		graph(8,6) <= "11111111";
		graph(8,7) <= "11111111";
		graph(8,8) <= "11111111";
		graph(8,9) <= "11111111";
		graph(8,10) <= "11111111";
		graph(8,11) <= "11111111";
		graph(8,12) <= "11111111";
		graph(8,13) <= "11111111";
		graph(8,14) <= "11111111";
		graph(8,15) <= "11111111";
		graph(8,16) <= "11111111";
		graph(8,17) <= "11111111";
		graph(8,18) <= "11111111";
		graph(8,19) <= "11111111";
		graph(8,20) <= "11111111";
		graph(8,21) <= "11111111";
		graph(8,22) <= "11111111";
		graph(8,23) <= "11111111";
		graph(8,24) <= "11111111";
		graph(8,25) <= "11111111";
		graph(8,26) <= "11111111";
		graph(8,27) <= "11111111";
		graph(8,28) <= "11111111";
		graph(8,29) <= "11111111";
		graph(8,30) <= "11111111";
		graph(8,31) <= "11111111";
		graph(9,0) <= "11111111";
		graph(9,1) <= "11111111";
		graph(9,2) <= "11111111";
		graph(9,3) <= "11111111";
		graph(9,4) <= "11111111";
		graph(9,5) <= "11111111";
		graph(9,6) <= "11111111";
		graph(9,7) <= "11111111";
		graph(9,8) <= "11111111";
		graph(9,9) <= "11111111";
		graph(9,10) <= "11111111";
		graph(9,11) <= "11111111";
		graph(9,12) <= "11111111";
		graph(9,13) <= "11111111";
		graph(9,14) <= "11111111";
		graph(9,15) <= "11111111";
		graph(9,16) <= "11111111";
		graph(9,17) <= "11111111";
		graph(9,18) <= "11111111";
		graph(9,19) <= "11111111";
		graph(9,20) <= "11111111";
		graph(9,21) <= "11111111";
		graph(9,22) <= "11111111";
		graph(9,23) <= "11111111";
		graph(9,24) <= "11111111";
		graph(9,25) <= "11111111";
		graph(9,26) <= "11111111";
		graph(9,27) <= "11111111";
		graph(9,28) <= "11111111";
		graph(9,29) <= "11111111";
		graph(9,30) <= "11111111";
		graph(9,31) <= "11111111";
		graph(10,0) <= "11111111";
		graph(10,1) <= "11111111";
		graph(10,2) <= "11111111";
		graph(10,3) <= "11111111";
		graph(10,4) <= "11111111";
		graph(10,5) <= "11111111";
		graph(10,6) <= "11111111";
		graph(10,7) <= "11111111";
		graph(10,8) <= "11111111";
		graph(10,9) <= "11111111";
		graph(10,10) <= "11111111";
		graph(10,11) <= "11111111";
		graph(10,12) <= "11111111";
		graph(10,13) <= "11111111";
		graph(10,14) <= "11111111";
		graph(10,15) <= "11111111";
		graph(10,16) <= "11111111";
		graph(10,17) <= "11111111";
		graph(10,18) <= "11111111";
		graph(10,19) <= "11111111";
		graph(10,20) <= "11111111";
		graph(10,21) <= "11111111";
		graph(10,22) <= "11111111";
		graph(10,23) <= "11111111";
		graph(10,24) <= "11111111";
		graph(10,25) <= "11111111";
		graph(10,26) <= "11111111";
		graph(10,27) <= "11111111";
		graph(10,28) <= "11111111";
		graph(10,29) <= "11111111";
		graph(10,30) <= "11111111";
		graph(10,31) <= "11111111";
		graph(11,0) <= "11111111";
		graph(11,1) <= "11111111";
		graph(11,2) <= "11111111";
		graph(11,3) <= "11111111";
		graph(11,4) <= "11111111";
		graph(11,5) <= "11111111";
		graph(11,6) <= "11111111";
		graph(11,7) <= "11111111";
		graph(11,8) <= "11111111";
		graph(11,9) <= "11111111";
		graph(11,10) <= "11111111";
		graph(11,11) <= "11111111";
		graph(11,12) <= "11111111";
		graph(11,13) <= "11111111";
		graph(11,14) <= "11111111";
		graph(11,15) <= "11111111";
		graph(11,16) <= "11111111";
		graph(11,17) <= "11111111";
		graph(11,18) <= "11111111";
		graph(11,19) <= "11111111";
		graph(11,20) <= "11111111";
		graph(11,21) <= "11111111";
		graph(11,22) <= "11111111";
		graph(11,23) <= "11111111";
		graph(11,24) <= "11111111";
		graph(11,25) <= "11111111";
		graph(11,26) <= "11111111";
		graph(11,27) <= "11111111";
		graph(11,28) <= "11111111";
		graph(11,29) <= "11111111";
		graph(11,30) <= "11111111";
		graph(11,31) <= "11111111";
		graph(12,0) <= "11111111";
		graph(12,1) <= "11111111";
		graph(12,2) <= "11111111";
		graph(12,3) <= "11111111";
		graph(12,4) <= "11111111";
		graph(12,5) <= "11111111";
		graph(12,6) <= "11111111";
		graph(12,7) <= "11111111";
		graph(12,8) <= "11111111";
		graph(12,9) <= "11111111";
		graph(12,10) <= "11111111";
		graph(12,11) <= "11111111";
		graph(12,12) <= "11111111";
		graph(12,13) <= "11111111";
		graph(12,14) <= "11111111";
		graph(12,15) <= "11111111";
		graph(12,16) <= "11111111";
		graph(12,17) <= "11111111";
		graph(12,18) <= "11111111";
		graph(12,19) <= "11111111";
		graph(12,20) <= "11111111";
		graph(12,21) <= "11111111";
		graph(12,22) <= "11111111";
		graph(12,23) <= "11111111";
		graph(12,24) <= "11111111";
		graph(12,25) <= "11111111";
		graph(12,26) <= "11111111";
		graph(12,27) <= "11111111";
		graph(12,28) <= "11111111";
		graph(12,29) <= "11111111";
		graph(12,30) <= "11111111";
		graph(12,31) <= "11111111";
		graph(13,0) <= "11111111";
		graph(13,1) <= "11111111";
		graph(13,2) <= "11111111";
		graph(13,3) <= "11111111";
		graph(13,4) <= "11111111";
		graph(13,5) <= "11111111";
		graph(13,6) <= "11111111";
		graph(13,7) <= "11111111";
		graph(13,8) <= "11111111";
		graph(13,9) <= "11111111";
		graph(13,10) <= "11111111";
		graph(13,11) <= "11111111";
		graph(13,12) <= "11111111";
		graph(13,13) <= "11111111";
		graph(13,14) <= "11111111";
		graph(13,15) <= "11111111";
		graph(13,16) <= "11111111";
		graph(13,17) <= "11111111";
		graph(13,18) <= "11111111";
		graph(13,19) <= "11111111";
		graph(13,20) <= "11111111";
		graph(13,21) <= "11111111";
		graph(13,22) <= "11111111";
		graph(13,23) <= "11111111";
		graph(13,24) <= "11111111";
		graph(13,25) <= "11111111";
		graph(13,26) <= "11111111";
		graph(13,27) <= "11111111";
		graph(13,28) <= "11111111";
		graph(13,29) <= "11111111";
		graph(13,30) <= "11111111";
		graph(13,31) <= "11111111";
		graph(14,0) <= "11111111";
		graph(14,1) <= "11111111";
		graph(14,2) <= "11111111";
		graph(14,3) <= "11111111";
		graph(14,4) <= "11111111";
		graph(14,5) <= "11111111";
		graph(14,6) <= "11111111";
		graph(14,7) <= "11111111";
		graph(14,8) <= "11111111";
		graph(14,9) <= "11111111";
		graph(14,10) <= "11111111";
		graph(14,11) <= "11111111";
		graph(14,12) <= "11111111";
		graph(14,13) <= "11111111";
		graph(14,14) <= "11111111";
		graph(14,15) <= "11111111";
		graph(14,16) <= "11111111";
		graph(14,17) <= "11111111";
		graph(14,18) <= "11111111";
		graph(14,19) <= "11111111";
		graph(14,20) <= "11111111";
		graph(14,21) <= "11111111";
		graph(14,22) <= "11111111";
		graph(14,23) <= "11111111";
		graph(14,24) <= "11111111";
		graph(14,25) <= "11111111";
		graph(14,26) <= "11111111";
		graph(14,27) <= "11111111";
		graph(14,28) <= "11111111";
		graph(14,29) <= "11111111";
		graph(14,30) <= "11111111";
		graph(14,31) <= "11111111";
		graph(15,0) <= "11111111";
		graph(15,1) <= "11111111";
		graph(15,2) <= "11111111";
		graph(15,3) <= "11111111";
		graph(15,4) <= "11111111";
		graph(15,5) <= "11111111";
		graph(15,6) <= "11111111";
		graph(15,7) <= "11111111";
		graph(15,8) <= "11111111";
		graph(15,9) <= "11111111";
		graph(15,10) <= "11111111";
		graph(15,11) <= "11111111";
		graph(15,12) <= "11111111";
		graph(15,13) <= "11111111";
		graph(15,14) <= "11111111";
		graph(15,15) <= "11111111";
		graph(15,16) <= "11111111";
		graph(15,17) <= "11111111";
		graph(15,18) <= "11111111";
		graph(15,19) <= "11111111";
		graph(15,20) <= "11111111";
		graph(15,21) <= "11111111";
		graph(15,22) <= "11111111";
		graph(15,23) <= "11111111";
		graph(15,24) <= "11111111";
		graph(15,25) <= "11111111";
		graph(15,26) <= "11111111";
		graph(15,27) <= "11111111";
		graph(15,28) <= "11111111";
		graph(15,29) <= "11111111";
		graph(15,30) <= "11111111";
		graph(15,31) <= "11111111";
		graph(16,0) <= "11111111";
		graph(16,1) <= "11111111";
		graph(16,2) <= "11111111";
		graph(16,3) <= "11111111";
		graph(16,4) <= "11111111";
		graph(16,5) <= "11111111";
		graph(16,6) <= "11111111";
		graph(16,7) <= "11111111";
		graph(16,8) <= "11111111";
		graph(16,9) <= "11111111";
		graph(16,10) <= "11111111";
		graph(16,11) <= "11111111";
		graph(16,12) <= "11111111";
		graph(16,13) <= "11111111";
		graph(16,14) <= "11111111";
		graph(16,15) <= "11111111";
		graph(16,16) <= "11111111";
		graph(16,17) <= "11111111";
		graph(16,18) <= "11111111";
		graph(16,19) <= "11111111";
		graph(16,20) <= "11111111";
		graph(16,21) <= "11111111";
		graph(16,22) <= "11111111";
		graph(16,23) <= "11111111";
		graph(16,24) <= "11111111";
		graph(16,25) <= "11111111";
		graph(16,26) <= "11111111";
		graph(16,27) <= "11111111";
		graph(16,28) <= "11111111";
		graph(16,29) <= "11111111";
		graph(16,30) <= "11111111";
		graph(16,31) <= "11111111";
		graph(17,0) <= "11111111";
		graph(17,1) <= "11111111";
		graph(17,2) <= "11111111";
		graph(17,3) <= "11111111";
		graph(17,4) <= "11111111";
		graph(17,5) <= "11111111";
		graph(17,6) <= "11111111";
		graph(17,7) <= "11111111";
		graph(17,8) <= "11111111";
		graph(17,9) <= "11111111";
		graph(17,10) <= "11111111";
		graph(17,11) <= "11111111";
		graph(17,12) <= "11111111";
		graph(17,13) <= "11111111";
		graph(17,14) <= "11111111";
		graph(17,15) <= "11111111";
		graph(17,16) <= "11111111";
		graph(17,17) <= "11111111";
		graph(17,18) <= "11111111";
		graph(17,19) <= "11111111";
		graph(17,20) <= "11111111";
		graph(17,21) <= "11111111";
		graph(17,22) <= "11111111";
		graph(17,23) <= "11111111";
		graph(17,24) <= "11111111";
		graph(17,25) <= "11111111";
		graph(17,26) <= "11111111";
		graph(17,27) <= "11111111";
		graph(17,28) <= "11111111";
		graph(17,29) <= "11111111";
		graph(17,30) <= "11111111";
		graph(17,31) <= "11111111";
		graph(18,0) <= "11111111";
		graph(18,1) <= "11111111";
		graph(18,2) <= "11111111";
		graph(18,3) <= "11111111";
		graph(18,4) <= "11111111";
		graph(18,5) <= "11111111";
		graph(18,6) <= "11111111";
		graph(18,7) <= "11111111";
		graph(18,8) <= "11111111";
		graph(18,9) <= "11111111";
		graph(18,10) <= "11111111";
		graph(18,11) <= "11111111";
		graph(18,12) <= "11111111";
		graph(18,13) <= "11111111";
		graph(18,14) <= "11111111";
		graph(18,15) <= "11111111";
		graph(18,16) <= "11111111";
		graph(18,17) <= "11111111";
		graph(18,18) <= "11111111";
		graph(18,19) <= "11111111";
		graph(18,20) <= "11111111";
		graph(18,21) <= "11111111";
		graph(18,22) <= "11111111";
		graph(18,23) <= "11111111";
		graph(18,24) <= "11111111";
		graph(18,25) <= "11111111";
		graph(18,26) <= "11111111";
		graph(18,27) <= "11111111";
		graph(18,28) <= "11111111";
		graph(18,29) <= "11111111";
		graph(18,30) <= "11111111";
		graph(18,31) <= "11111111";
		graph(19,0) <= "11111111";
		graph(19,1) <= "11111111";
		graph(19,2) <= "11111111";
		graph(19,3) <= "11111111";
		graph(19,4) <= "11111111";
		graph(19,5) <= "11111111";
		graph(19,6) <= "11111111";
		graph(19,7) <= "11111111";
		graph(19,8) <= "11111111";
		graph(19,9) <= "11111111";
		graph(19,10) <= "11111111";
		graph(19,11) <= "11111111";
		graph(19,12) <= "11111111";
		graph(19,13) <= "11111111";
		graph(19,14) <= "11111111";
		graph(19,15) <= "11111111";
		graph(19,16) <= "11111111";
		graph(19,17) <= "11111111";
		graph(19,18) <= "11111111";
		graph(19,19) <= "11111111";
		graph(19,20) <= "11111111";
		graph(19,21) <= "11111111";
		graph(19,22) <= "11111111";
		graph(19,23) <= "11111111";
		graph(19,24) <= "11111111";
		graph(19,25) <= "11111111";
		graph(19,26) <= "11111111";
		graph(19,27) <= "11111111";
		graph(19,28) <= "11111111";
		graph(19,29) <= "11111111";
		graph(19,30) <= "11111111";
		graph(19,31) <= "11111111";
		graph(20,0) <= "11111111";
		graph(20,1) <= "11111111";
		graph(20,2) <= "11111111";
		graph(20,3) <= "11111111";
		graph(20,4) <= "11111111";
		graph(20,5) <= "11111111";
		graph(20,6) <= "11111111";
		graph(20,7) <= "11111111";
		graph(20,8) <= "11111111";
		graph(20,9) <= "11111111";
		graph(20,10) <= "11111111";
		graph(20,11) <= "11111111";
		graph(20,12) <= "11111111";
		graph(20,13) <= "11111111";
		graph(20,14) <= "11111111";
		graph(20,15) <= "11111111";
		graph(20,16) <= "11111111";
		graph(20,17) <= "11111111";
		graph(20,18) <= "11111111";
		graph(20,19) <= "11111111";
		graph(20,20) <= "11111111";
		graph(20,21) <= "11111111";
		graph(20,22) <= "11111111";
		graph(20,23) <= "11111111";
		graph(20,24) <= "11111111";
		graph(20,25) <= "11111111";
		graph(20,26) <= "11111111";
		graph(20,27) <= "11111111";
		graph(20,28) <= "11111111";
		graph(20,29) <= "11111111";
		graph(20,30) <= "11111111";
		graph(20,31) <= "11111111";
		graph(21,0) <= "11111111";
		graph(21,1) <= "11111111";
		graph(21,2) <= "11111111";
		graph(21,3) <= "11111111";
		graph(21,4) <= "11111111";
		graph(21,5) <= "11111111";
		graph(21,6) <= "11111111";
		graph(21,7) <= "11111111";
		graph(21,8) <= "11111111";
		graph(21,9) <= "11111111";
		graph(21,10) <= "11111111";
		graph(21,11) <= "11111111";
		graph(21,12) <= "11111111";
		graph(21,13) <= "11111111";
		graph(21,14) <= "11111111";
		graph(21,15) <= "11111111";
		graph(21,16) <= "11111111";
		graph(21,17) <= "11111111";
		graph(21,18) <= "11111111";
		graph(21,19) <= "11111111";
		graph(21,20) <= "11111111";
		graph(21,21) <= "11111111";
		graph(21,22) <= "11111111";
		graph(21,23) <= "11111111";
		graph(21,24) <= "11111111";
		graph(21,25) <= "11111111";
		graph(21,26) <= "11111111";
		graph(21,27) <= "11111111";
		graph(21,28) <= "11111111";
		graph(21,29) <= "11111111";
		graph(21,30) <= "11111111";
		graph(21,31) <= "11111111";
		graph(22,0) <= "11111111";
		graph(22,1) <= "11111111";
		graph(22,2) <= "11111111";
		graph(22,3) <= "11111111";
		graph(22,4) <= "11111111";
		graph(22,5) <= "11111111";
		graph(22,6) <= "11111111";
		graph(22,7) <= "11111111";
		graph(22,8) <= "11111111";
		graph(22,9) <= "11111111";
		graph(22,10) <= "11111111";
		graph(22,11) <= "11111111";
		graph(22,12) <= "11111111";
		graph(22,13) <= "11111111";
		graph(22,14) <= "11111111";
		graph(22,15) <= "11111111";
		graph(22,16) <= "11111111";
		graph(22,17) <= "11111111";
		graph(22,18) <= "11111111";
		graph(22,19) <= "11111111";
		graph(22,20) <= "11111111";
		graph(22,21) <= "11111111";
		graph(22,22) <= "11111111";
		graph(22,23) <= "11111111";
		graph(22,24) <= "11111111";
		graph(22,25) <= "11111111";
		graph(22,26) <= "11111111";
		graph(22,27) <= "11111111";
		graph(22,28) <= "11111111";
		graph(22,29) <= "11111111";
		graph(22,30) <= "11111111";
		graph(22,31) <= "11111111";
		graph(23,0) <= "11111111";
		graph(23,1) <= "11111111";
		graph(23,2) <= "11111111";
		graph(23,3) <= "11111111";
		graph(23,4) <= "11111111";
		graph(23,5) <= "11111111";
		graph(23,6) <= "11111111";
		graph(23,7) <= "11111111";
		graph(23,8) <= "11111111";
		graph(23,9) <= "11111111";
		graph(23,10) <= "11111111";
		graph(23,11) <= "11111111";
		graph(23,12) <= "11111111";
		graph(23,13) <= "11111111";
		graph(23,14) <= "11111111";
		graph(23,15) <= "11111111";
		graph(23,16) <= "11111111";
		graph(23,17) <= "11111111";
		graph(23,18) <= "11111111";
		graph(23,19) <= "11111111";
		graph(23,20) <= "11111111";
		graph(23,21) <= "11111111";
		graph(23,22) <= "11111111";
		graph(23,23) <= "11111111";
		graph(23,24) <= "11111111";
		graph(23,25) <= "11111111";
		graph(23,26) <= "11111111";
		graph(23,27) <= "11111111";
		graph(23,28) <= "11111111";
		graph(23,29) <= "11111111";
		graph(23,30) <= "11111111";
		graph(23,31) <= "11111111";
		graph(24,0) <= "11111111";
		graph(24,1) <= "11111111";
		graph(24,2) <= "11111111";
		graph(24,3) <= "11111111";
		graph(24,4) <= "11111111";
		graph(24,5) <= "11111111";
		graph(24,6) <= "11111111";
		graph(24,7) <= "11111111";
		graph(24,8) <= "11111111";
		graph(24,9) <= "11111111";
		graph(24,10) <= "11111111";
		graph(24,11) <= "11111111";
		graph(24,12) <= "11111111";
		graph(24,13) <= "11111111";
		graph(24,14) <= "11111111";
		graph(24,15) <= "11111111";
		graph(24,16) <= "11111111";
		graph(24,17) <= "11111111";
		graph(24,18) <= "11111111";
		graph(24,19) <= "11111111";
		graph(24,20) <= "11111111";
		graph(24,21) <= "11111111";
		graph(24,22) <= "11111111";
		graph(24,23) <= "11111111";
		graph(24,24) <= "11111111";
		graph(24,25) <= "11111111";
		graph(24,26) <= "11111111";
		graph(24,27) <= "11111111";
		graph(24,28) <= "11111111";
		graph(24,29) <= "11111111";
		graph(24,30) <= "11111111";
		graph(24,31) <= "11111111";
		graph(25,0) <= "11111111";
		graph(25,1) <= "11111111";
		graph(25,2) <= "11111111";
		graph(25,3) <= "11111111";
		graph(25,4) <= "11111111";
		graph(25,5) <= "11111111";
		graph(25,6) <= "11111111";
		graph(25,7) <= "11111111";
		graph(25,8) <= "11111111";
		graph(25,9) <= "11111111";
		graph(25,10) <= "11111111";
		graph(25,11) <= "11111111";
		graph(25,12) <= "11111111";
		graph(25,13) <= "11111111";
		graph(25,14) <= "11111111";
		graph(25,15) <= "11111111";
		graph(25,16) <= "11111111";
		graph(25,17) <= "11111111";
		graph(25,18) <= "11111111";
		graph(25,19) <= "11111111";
		graph(25,20) <= "11111111";
		graph(25,21) <= "11111111";
		graph(25,22) <= "11111111";
		graph(25,23) <= "11111111";
		graph(25,24) <= "11111111";
		graph(25,25) <= "11111111";
		graph(25,26) <= "11111111";
		graph(25,27) <= "11111111";
		graph(25,28) <= "11111111";
		graph(25,29) <= "11111111";
		graph(25,30) <= "11111111";
		graph(25,31) <= "11111111";
		graph(26,0) <= "11111111";
		graph(26,1) <= "11111111";
		graph(26,2) <= "11111111";
		graph(26,3) <= "11111111";
		graph(26,4) <= "11111111";
		graph(26,5) <= "11111111";
		graph(26,6) <= "11111111";
		graph(26,7) <= "11111111";
		graph(26,8) <= "11111111";
		graph(26,9) <= "11111111";
		graph(26,10) <= "11111111";
		graph(26,11) <= "11111111";
		graph(26,12) <= "11111111";
		graph(26,13) <= "11111111";
		graph(26,14) <= "11111111";
		graph(26,15) <= "11111111";
		graph(26,16) <= "11111111";
		graph(26,17) <= "11111111";
		graph(26,18) <= "11111111";
		graph(26,19) <= "11111111";
		graph(26,20) <= "11111111";
		graph(26,21) <= "11111111";
		graph(26,22) <= "11111111";
		graph(26,23) <= "11111111";
		graph(26,24) <= "11111111";
		graph(26,25) <= "11111111";
		graph(26,26) <= "11111111";
		graph(26,27) <= "11111111";
		graph(26,28) <= "11111111";
		graph(26,29) <= "11111111";
		graph(26,30) <= "11111111";
		graph(26,31) <= "11111111";
		graph(27,0) <= "11111111";
		graph(27,1) <= "11111111";
		graph(27,2) <= "11111111";
		graph(27,3) <= "11111111";
		graph(27,4) <= "11111111";
		graph(27,5) <= "11111111";
		graph(27,6) <= "11111111";
		graph(27,7) <= "11111111";
		graph(27,8) <= "11111111";
		graph(27,9) <= "11111111";
		graph(27,10) <= "11111111";
		graph(27,11) <= "11111111";
		graph(27,12) <= "11111111";
		graph(27,13) <= "11111111";
		graph(27,14) <= "11111111";
		graph(27,15) <= "11111111";
		graph(27,16) <= "11111111";
		graph(27,17) <= "11111111";
		graph(27,18) <= "11111111";
		graph(27,19) <= "11111111";
		graph(27,20) <= "11111111";
		graph(27,21) <= "11111111";
		graph(27,22) <= "11111111";
		graph(27,23) <= "11111111";
		graph(27,24) <= "11111111";
		graph(27,25) <= "11111111";
		graph(27,26) <= "11111111";
		graph(27,27) <= "11111111";
		graph(27,28) <= "11111111";
		graph(27,29) <= "11111111";
		graph(27,30) <= "11111111";
		graph(27,31) <= "11111111";
		graph(28,0) <= "11111111";
		graph(28,1) <= "11111111";
		graph(28,2) <= "11111111";
		graph(28,3) <= "11111111";
		graph(28,4) <= "11111111";
		graph(28,5) <= "11111111";
		graph(28,6) <= "11111111";
		graph(28,7) <= "11111111";
		graph(28,8) <= "11111111";
		graph(28,9) <= "11111111";
		graph(28,10) <= "11111111";
		graph(28,11) <= "11111111";
		graph(28,12) <= "11111111";
		graph(28,13) <= "11111111";
		graph(28,14) <= "11111111";
		graph(28,15) <= "11111111";
		graph(28,16) <= "11111111";
		graph(28,17) <= "11111111";
		graph(28,18) <= "11111111";
		graph(28,19) <= "11111111";
		graph(28,20) <= "11111111";
		graph(28,21) <= "11111111";
		graph(28,22) <= "11111111";
		graph(28,23) <= "11111111";
		graph(28,24) <= "11111111";
		graph(28,25) <= "11111111";
		graph(28,26) <= "11111111";
		graph(28,27) <= "11111111";
		graph(28,28) <= "11111111";
		graph(28,29) <= "11111111";
		graph(28,30) <= "11111111";
		graph(28,31) <= "11111111";
		graph(29,0) <= "11111111";
		graph(29,1) <= "11111111";
		graph(29,2) <= "11111111";
		graph(29,3) <= "11111111";
		graph(29,4) <= "11111111";
		graph(29,5) <= "11111111";
		graph(29,6) <= "11111111";
		graph(29,7) <= "11111111";
		graph(29,8) <= "11111111";
		graph(29,9) <= "11111111";
		graph(29,10) <= "11111111";
		graph(29,11) <= "11111111";
		graph(29,12) <= "11111111";
		graph(29,13) <= "11111111";
		graph(29,14) <= "11111111";
		graph(29,15) <= "11111111";
		graph(29,16) <= "11111111";
		graph(29,17) <= "11111111";
		graph(29,18) <= "11111111";
		graph(29,19) <= "11111111";
		graph(29,20) <= "11111111";
		graph(29,21) <= "11111111";
		graph(29,22) <= "11111111";
		graph(29,23) <= "11111111";
		graph(29,24) <= "11111111";
		graph(29,25) <= "11111111";
		graph(29,26) <= "11111111";
		graph(29,27) <= "11111111";
		graph(29,28) <= "11111111";
		graph(29,29) <= "11111111";
		graph(29,30) <= "11111111";
		graph(29,31) <= "11111111";
		graph(30,0) <= "11111111";
		graph(30,1) <= "11111111";
		graph(30,2) <= "11111111";
		graph(30,3) <= "11111111";
		graph(30,4) <= "11111111";
		graph(30,5) <= "11111111";
		graph(30,6) <= "11111111";
		graph(30,7) <= "11111111";
		graph(30,8) <= "11111111";
		graph(30,9) <= "11111111";
		graph(30,10) <= "11111111";
		graph(30,11) <= "11111111";
		graph(30,12) <= "11111111";
		graph(30,13) <= "11111111";
		graph(30,14) <= "11111111";
		graph(30,15) <= "11111111";
		graph(30,16) <= "11111111";
		graph(30,17) <= "11111111";
		graph(30,18) <= "11111111";
		graph(30,19) <= "11111111";
		graph(30,20) <= "11111111";
		graph(30,21) <= "11111111";
		graph(30,22) <= "11111111";
		graph(30,23) <= "11111111";
		graph(30,24) <= "11111111";
		graph(30,25) <= "11111111";
		graph(30,26) <= "11111111";
		graph(30,27) <= "11111111";
		graph(30,28) <= "11111111";
		graph(30,29) <= "11111111";
		graph(30,30) <= "11111111";
		graph(30,31) <= "11111111";
		graph(31,0) <= "11111111";
		graph(31,1) <= "11111111";
		graph(31,2) <= "11111111";
		graph(31,3) <= "11111111";
		graph(31,4) <= "11111111";
		graph(31,5) <= "11111111";
		graph(31,6) <= "11111111";
		graph(31,7) <= "11111111";
		graph(31,8) <= "11111111";
		graph(31,9) <= "11111111";
		graph(31,10) <= "11111111";
		graph(31,11) <= "11111111";
		graph(31,12) <= "11111111";
		graph(31,13) <= "11111111";
		graph(31,14) <= "11111111";
		graph(31,15) <= "11111111";
		graph(31,16) <= "11111111";
		graph(31,17) <= "11111111";
		graph(31,18) <= "11111111";
		graph(31,19) <= "11111111";
		graph(31,20) <= "11111111";
		graph(31,21) <= "11111111";
		graph(31,22) <= "11111111";
		graph(31,23) <= "11111111";
		graph(31,24) <= "11111111";
		graph(31,25) <= "11111111";
		graph(31,26) <= "11111111";
		graph(31,27) <= "11111111";
		graph(31,28) <= "11111111";
		graph(31,29) <= "11111111";
		graph(31,30) <= "11111111";
		graph(31,31) <= "11111111";

		d1 := DD(0, 4);
		d2 := DD(0, 5);
		d3 := DD(0, 6);
		d4 := DD(0, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(0, 0);
		e2 := DD(0, 1);
		e3 := DD(0, 2);
		e4 := DD(0, 3);
		e := e1 & e2 & e3 & e4;

		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(1, 4);
		d2 := DD(1, 5);
		d3 := DD(1, 6); 
		d4 := DD(1, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(1, 0);
		e2 := DD(1, 1);
		e3 := DD(1, 2);
		e4 := DD(1, 3);
		e := e1 & e2 & e3 & e4;
		
		--report "here1";
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(2, 4);
		d2 := DD(2, 5);
		d3 := DD(2, 6);
		d4 := DD(2, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(2, 0);
		e2 := DD(2, 1);
		e3 := DD(2, 2);
		e4 := DD(2, 3);
		e := e1 & e2 & e3 & e4;
		
		--report "here2";
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(3, 4);
		d2 := DD(3, 5);
		d3 := DD(3, 6);
		d4 := DD(3, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(3, 0);
		e2 := DD(3, 1);
		e3 := DD(3, 2);
		e4 := DD(3, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(4, 4);
		d2 := DD(4, 5);
		d3 := DD(4, 6);
		d4 := DD(4, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(4, 0);
		e2 := DD(4, 1);
		e3 := DD(4, 2);
		e4 := DD(4, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(5, 4);
		d2 := DD(5, 5);
		d3 := DD(5, 6);
		d4 := DD(5, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(5, 0);
		e2 := DD(5, 1);
		e3 := DD(5, 2);
		e4 := DD(5, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(6, 4);
		d2 := DD(6, 5);
		d3 := DD(6, 6);
		d4 := DD(6, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(6, 0);
		e2 := DD(6, 1);
		e3 := DD(6, 2);
		e4 := DD(6, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(7, 4);
		d2 := DD(7, 5);
		d3 := DD(7, 6);
		d4 := DD(7, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(7, 0);
		e2 := DD(7, 1);
		e3 := DD(7, 2);
		e4 := DD(7, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(8, 4);
		d2 := DD(8, 5);
		d3 := DD(8, 6);
		d4 := DD(8, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(8, 0);
		e2 := DD(8, 1);
		e3 := DD(8, 2);
		e4 := DD(8, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(9, 4);
		d2 := DD(9, 5);
		d3 := DD(9, 6);
		d4 := DD(9, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(9, 0);
		e2 := DD(9, 1);
		e3 := DD(9, 2);
		e4 := DD(9, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(10, 4);
		d2 := DD(10, 5);
		d3 := DD(10, 6);
		d4 := DD(10, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(10, 0);
		e2 := DD(10, 1);
		e3 := DD(10, 2);
		e4 := DD(10, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(11, 4);
		d2 := DD(11, 5);
		d3 := DD(11, 6);
		d4 := DD(11, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(11, 0);
		e2 := DD(11, 1);
		e3 := DD(11, 2);
		e4 := DD(11, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(12, 4);
		d2 := DD(12, 5);
		d3 := DD(12, 6);
		d4 := DD(12, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(12, 0);
		e2 := DD(12, 1);
		e3 := DD(12, 2);
		e4 := DD(12, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(13, 4);
		d2 := DD(13, 5);
		d3 := DD(13, 6);
		d4 := DD(13, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(13, 0);
		e2 := DD(13, 1);
		e3 := DD(13, 2);
		e4 := DD(13, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(14, 4);
		d2 := DD(14, 5);
		d3 := DD(14, 6);
		d4 := DD(14, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(14, 0);
		e2 := DD(14, 1);
		e3 := DD(14, 2);
		e4 := DD(14, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(15, 4);
		d2 := DD(15, 5);
		d3 := DD(15, 6);
		d4 := DD(15, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(15, 0);
		e2 := DD(15, 1);
		e3 := DD(15, 2);
		e4 := DD(15, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(16, 4);
		d2 := DD(16, 5);
		d3 := DD(16, 6);
		d4 := DD(16, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(16, 0);
		e2 := DD(16, 1);
		e3 := DD(16, 2);
		e4 := DD(16, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(17, 4);
		d2 := DD(17, 5);
		d3 := DD(17, 6);
		d4 := DD(17, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(17, 0);
		e2 := DD(17, 1);
		e3 := DD(17, 2);
		e4 := DD(17, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(18, 4);
		d2 := DD(18, 5);
		d3 := DD(18, 6);
		d4 := DD(18, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(18, 0);
		e2 := DD(18, 1);
		e3 := DD(18, 2);
		e4 := DD(18, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(19, 4);
		d2 := DD(19, 5);
		d3 := DD(19, 6);
		d4 := DD(19, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(19, 0);
		e2 := DD(19, 1);
		e3 := DD(19, 2);
		e4 := DD(19, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(20, 4);
		d2 := DD(20, 5);
		d3 := DD(20, 6);
		d4 := DD(20, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(20, 0);
		e2 := DD(20, 1);
		e3 := DD(20, 2);
		e4 := DD(20, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(21, 4);
		d2 := DD(21, 5);
		d3 := DD(21, 6);
		d4 := DD(21, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(21, 0);
		e2 := DD(21, 1);
		e3 := DD(21, 2);
		e4 := DD(21, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(22, 4);
		d2 := DD(22, 5);
		d3 := DD(22, 6);
		d4 := DD(22, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(22, 0);
		e2 := DD(22, 1);
		e3 := DD(22, 2);
		e4 := DD(22, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(23, 4);
		d2 := DD(23, 5);
		d3 := DD(23, 6);
		d4 := DD(23, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(23, 0);
		e2 := DD(23, 1);
		e3 := DD(23, 2);
		e4 := DD(23, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(24, 4);
		d2 := DD(24, 5);
		d3 := DD(24, 6);
		d4 := DD(24, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(24, 0);
		e2 := DD(24, 1);
		e3 := DD(24, 2);
		e4 := DD(24, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(25, 4);
		d2 := DD(25, 5);
		d3 := DD(25, 6);
		d4 := DD(25, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(25, 0);
		e2 := DD(25, 1);
		e3 := DD(25, 2);
		e4 := DD(25, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(26, 4);
		d2 := DD(26, 5);
		d3 := DD(26, 6);
		d4 := DD(26, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(26, 0);
		e2 := DD(26, 1);
		e3 := DD(26, 2);
		e4 := DD(26, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(27, 4);
		d2 := DD(27, 5);
		d3 := DD(27, 6);
		d4 := DD(27, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(27, 0);
		e2 := DD(27, 1);
		e3 := DD(27, 2);
		e4 := DD(27, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(28, 4);
		d2 := DD(28, 5);
		d3 := DD(28, 6);
		d4 := DD(28, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(28, 0);
		e2 := DD(28, 1);
		e3 := DD(28, 2);
		e4 := DD(28, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(29, 4);
		d2 := DD(29, 5);
		d3 := DD(29, 6);
		d4 := DD(29, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(29, 0);
		e2 := DD(29, 1);
		e3 := DD(29, 2);
		e4 := DD(29, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(30, 4);
		d2 := DD(30, 5);
		d3 := DD(30, 6);
		d4 := DD(30, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(30, 0);
		e2 := DD(30, 1);
		e3 := DD(30, 2);
		e4 := DD(30, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;
		d1 := DD(31, 4);
		d2 := DD(31, 5);
		d3 := DD(31, 6);
		d4 := DD(31, 7);
		d := d1 & d2 & d3 & d4;
		e1 := DD(31, 0);
		e2 := DD(31, 1);
		e3 := DD(31, 2);
		e4 := DD(31, 3);
		e := e1 & e2 & e3 & e4;
		IP_ADDR(to_integer(unsigned(d))) <= e;

		-- Manipulating graph entries

		d1 := DD(0, 12);
		d2 := DD(0, 13);
		d3 := DD(0, 14);
		d4 := DD(0, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 21);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(0, 22);
		d2 := DD(0, 23);
		d3 := DD(0, 24);
		d4 := DD(0, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 31);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(0, 32);
		d2 := DD(0, 33);
		d3 := DD(0, 34);
		d4 := DD(0, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 41);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(0, 42);
		d2 := DD(0, 43);
		d3 := DD(0, 44);
		d4 := DD(0, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 51);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(0, 52);
		d2 := DD(0, 53);
		d3 := DD(0, 54);
		d4 := DD(0, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 61);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(0, 62);
		d2 := DD(0, 63);
		d3 := DD(0, 64);
		d4 := DD(0, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 71);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(0, 72);
		d2 := DD(0, 73);
		d3 := DD(0, 74);
		d4 := DD(0, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 81);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(0, 82);
		d2 := DD(0, 83);
		d3 := DD(0, 84);
		d4 := DD(0, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(0, 91);
		graph(0, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 12);
		d2 := DD(1, 13);
		d3 := DD(1, 14);
		d4 := DD(1, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 21);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 22);
		d2 := DD(1, 23);
		d3 := DD(1, 24);
		d4 := DD(1, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 31);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 32);
		d2 := DD(1, 33);
		d3 := DD(1, 34);
		d4 := DD(1, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 41);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 42);
		d2 := DD(1, 43);
		d3 := DD(1, 44);
		d4 := DD(1, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 51);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 52);
		d2 := DD(1, 53);
		d3 := DD(1, 54);
		d4 := DD(1, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 61);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 62);
		d2 := DD(1, 63);
		d3 := DD(1, 64);
		d4 := DD(1, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 71);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 72);
		d2 := DD(1, 73);
		d3 := DD(1, 74);
		d4 := DD(1, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 81);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(1, 82);
		d2 := DD(1, 83);
		d3 := DD(1, 84);
		d4 := DD(1, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(1, 91);
		graph(1, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 12);
		d2 := DD(2, 13);
		d3 := DD(2, 14);
		d4 := DD(2, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 21);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 22);
		d2 := DD(2, 23);
		d3 := DD(2, 24);
		d4 := DD(2, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 31);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 32);
		d2 := DD(2, 33);
		d3 := DD(2, 34);
		d4 := DD(2, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 41);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 42);
		d2 := DD(2, 43);
		d3 := DD(2, 44);
		d4 := DD(2, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 51);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 52);
		d2 := DD(2, 53);
		d3 := DD(2, 54);
		d4 := DD(2, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 61);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 62);
		d2 := DD(2, 63);
		d3 := DD(2, 64);
		d4 := DD(2, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 71);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 72);
		d2 := DD(2, 73);
		d3 := DD(2, 74);
		d4 := DD(2, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 81);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(2, 82);
		d2 := DD(2, 83);
		d3 := DD(2, 84);
		d4 := DD(2, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(2, 91);
		graph(2, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 12);
		d2 := DD(3, 13);
		d3 := DD(3, 14);
		d4 := DD(3, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 21);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 22);
		d2 := DD(3, 23);
		d3 := DD(3, 24);
		d4 := DD(3, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 31);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 32);
		d2 := DD(3, 33);
		d3 := DD(3, 34);
		d4 := DD(3, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 41);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 42);
		d2 := DD(3, 43);
		d3 := DD(3, 44);
		d4 := DD(3, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 51);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 52);
		d2 := DD(3, 53);
		d3 := DD(3, 54);
		d4 := DD(3, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 61);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 62);
		d2 := DD(3, 63);
		d3 := DD(3, 64);
		d4 := DD(3, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 71);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 72);
		d2 := DD(3, 73);
		d3 := DD(3, 74);
		d4 := DD(3, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 81);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(3, 82);
		d2 := DD(3, 83);
		d3 := DD(3, 84);
		d4 := DD(3, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(3, 91);
		graph(3, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 12);
		d2 := DD(4, 13);
		d3 := DD(4, 14);
		d4 := DD(4, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 21);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 22);
		d2 := DD(4, 23);
		d3 := DD(4, 24);
		d4 := DD(4, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 31);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 32);
		d2 := DD(4, 33);
		d3 := DD(4, 34);
		d4 := DD(4, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 41);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 42);
		d2 := DD(4, 43);
		d3 := DD(4, 44);
		d4 := DD(4, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 51);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 52);
		d2 := DD(4, 53);
		d3 := DD(4, 54);
		d4 := DD(4, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 61);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 62);
		d2 := DD(4, 63);
		d3 := DD(4, 64);
		d4 := DD(4, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 71);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 72);
		d2 := DD(4, 73);
		d3 := DD(4, 74);
		d4 := DD(4, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 81);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(4, 82);
		d2 := DD(4, 83);
		d3 := DD(4, 84);
		d4 := DD(4, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(4, 91);
		graph(4, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 12);
		d2 := DD(5, 13);
		d3 := DD(5, 14);
		d4 := DD(5, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 21);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 22);
		d2 := DD(5, 23);
		d3 := DD(5, 24);
		d4 := DD(5, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 31);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 32);
		d2 := DD(5, 33);
		d3 := DD(5, 34);
		d4 := DD(5, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 41);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 42);
		d2 := DD(5, 43);
		d3 := DD(5, 44);
		d4 := DD(5, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 51);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 52);
		d2 := DD(5, 53);
		d3 := DD(5, 54);
		d4 := DD(5, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 61);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 62);
		d2 := DD(5, 63);
		d3 := DD(5, 64);
		d4 := DD(5, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 71);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 72);
		d2 := DD(5, 73);
		d3 := DD(5, 74);
		d4 := DD(5, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 81);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(5, 82);
		d2 := DD(5, 83);
		d3 := DD(5, 84);
		d4 := DD(5, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(5, 91);
		graph(5, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 12);
		d2 := DD(6, 13);
		d3 := DD(6, 14);
		d4 := DD(6, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 21);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 22);
		d2 := DD(6, 23);
		d3 := DD(6, 24);
		d4 := DD(6, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 31);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 32);
		d2 := DD(6, 33);
		d3 := DD(6, 34);
		d4 := DD(6, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 41);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 42);
		d2 := DD(6, 43);
		d3 := DD(6, 44);
		d4 := DD(6, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 51);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 52);
		d2 := DD(6, 53);
		d3 := DD(6, 54);
		d4 := DD(6, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 61);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 62);
		d2 := DD(6, 63);
		d3 := DD(6, 64);
		d4 := DD(6, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 71);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 72);
		d2 := DD(6, 73);
		d3 := DD(6, 74);
		d4 := DD(6, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 81);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(6, 82);
		d2 := DD(6, 83);
		d3 := DD(6, 84);
		d4 := DD(6, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(6, 91);
		graph(6, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 12);
		d2 := DD(7, 13);
		d3 := DD(7, 14);
		d4 := DD(7, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 21);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 22);
		d2 := DD(7, 23);
		d3 := DD(7, 24);
		d4 := DD(7, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 31);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 32);
		d2 := DD(7, 33);
		d3 := DD(7, 34);
		d4 := DD(7, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 41);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 42);
		d2 := DD(7, 43);
		d3 := DD(7, 44);
		d4 := DD(7, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 51);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 52);
		d2 := DD(7, 53);
		d3 := DD(7, 54);
		d4 := DD(7, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 61);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 62);
		d2 := DD(7, 63);
		d3 := DD(7, 64);
		d4 := DD(7, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 71);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 72);
		d2 := DD(7, 73);
		d3 := DD(7, 74);
		d4 := DD(7, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 81);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(7, 82);
		d2 := DD(7, 83);
		d3 := DD(7, 84);
		d4 := DD(7, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(7, 91);
		graph(7, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 12);
		d2 := DD(8, 13);
		d3 := DD(8, 14);
		d4 := DD(8, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 21);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 22);
		d2 := DD(8, 23);
		d3 := DD(8, 24);
		d4 := DD(8, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 31);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 32);
		d2 := DD(8, 33);
		d3 := DD(8, 34);
		d4 := DD(8, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 41);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 42);
		d2 := DD(8, 43);
		d3 := DD(8, 44);
		d4 := DD(8, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 51);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 52);
		d2 := DD(8, 53);
		d3 := DD(8, 54);
		d4 := DD(8, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 61);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 62);
		d2 := DD(8, 63);
		d3 := DD(8, 64);
		d4 := DD(8, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 71);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 72);
		d2 := DD(8, 73);
		d3 := DD(8, 74);
		d4 := DD(8, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 81);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(8, 82);
		d2 := DD(8, 83);
		d3 := DD(8, 84);
		d4 := DD(8, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(8, 91);
		graph(8, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 12);
		d2 := DD(9, 13);
		d3 := DD(9, 14);
		d4 := DD(9, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 21);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 22);
		d2 := DD(9, 23);
		d3 := DD(9, 24);
		d4 := DD(9, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 31);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 32);
		d2 := DD(9, 33);
		d3 := DD(9, 34);
		d4 := DD(9, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 41);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 42);
		d2 := DD(9, 43);
		d3 := DD(9, 44);
		d4 := DD(9, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 51);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 52);
		d2 := DD(9, 53);
		d3 := DD(9, 54);
		d4 := DD(9, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 61);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 62);
		d2 := DD(9, 63);
		d3 := DD(9, 64);
		d4 := DD(9, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 71);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 72);
		d2 := DD(9, 73);
		d3 := DD(9, 74);
		d4 := DD(9, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 81);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(9, 82);
		d2 := DD(9, 83);
		d3 := DD(9, 84);
		d4 := DD(9, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(9, 91);
		graph(9, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 12);
		d2 := DD(10, 13);
		d3 := DD(10, 14);
		d4 := DD(10, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 21);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 22);
		d2 := DD(10, 23);
		d3 := DD(10, 24);
		d4 := DD(10, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 31);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 32);
		d2 := DD(10, 33);
		d3 := DD(10, 34);
		d4 := DD(10, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 41);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 42);
		d2 := DD(10, 43);
		d3 := DD(10, 44);
		d4 := DD(10, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 51);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 52);
		d2 := DD(10, 53);
		d3 := DD(10, 54);
		d4 := DD(10, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 61);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 62);
		d2 := DD(10, 63);
		d3 := DD(10, 64);
		d4 := DD(10, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 71);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 72);
		d2 := DD(10, 73);
		d3 := DD(10, 74);
		d4 := DD(10, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 81);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(10, 82);
		d2 := DD(10, 83);
		d3 := DD(10, 84);
		d4 := DD(10, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(10, 91);
		graph(10, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 12);
		d2 := DD(11, 13);
		d3 := DD(11, 14);
		d4 := DD(11, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 21);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 22);
		d2 := DD(11, 23);
		d3 := DD(11, 24);
		d4 := DD(11, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 31);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 32);
		d2 := DD(11, 33);
		d3 := DD(11, 34);
		d4 := DD(11, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 41);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 42);
		d2 := DD(11, 43);
		d3 := DD(11, 44);
		d4 := DD(11, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 51);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 52);
		d2 := DD(11, 53);
		d3 := DD(11, 54);
		d4 := DD(11, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 61);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 62);
		d2 := DD(11, 63);
		d3 := DD(11, 64);
		d4 := DD(11, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 71);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 72);
		d2 := DD(11, 73);
		d3 := DD(11, 74);
		d4 := DD(11, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 81);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(11, 82);
		d2 := DD(11, 83);
		d3 := DD(11, 84);
		d4 := DD(11, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(11, 91);
		graph(11, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 12);
		d2 := DD(12, 13);
		d3 := DD(12, 14);
		d4 := DD(12, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 21);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 22);
		d2 := DD(12, 23);
		d3 := DD(12, 24);
		d4 := DD(12, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 31);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 32);
		d2 := DD(12, 33);
		d3 := DD(12, 34);
		d4 := DD(12, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 41);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 42);
		d2 := DD(12, 43);
		d3 := DD(12, 44);
		d4 := DD(12, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 51);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 52);
		d2 := DD(12, 53);
		d3 := DD(12, 54);
		d4 := DD(12, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 61);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 62);
		d2 := DD(12, 63);
		d3 := DD(12, 64);
		d4 := DD(12, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 71);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 72);
		d2 := DD(12, 73);
		d3 := DD(12, 74);
		d4 := DD(12, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 81);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(12, 82);
		d2 := DD(12, 83);
		d3 := DD(12, 84);
		d4 := DD(12, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(12, 91);
		graph(12, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 12);
		d2 := DD(13, 13);
		d3 := DD(13, 14);
		d4 := DD(13, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 21);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 22);
		d2 := DD(13, 23);
		d3 := DD(13, 24);
		d4 := DD(13, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 31);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 32);
		d2 := DD(13, 33);
		d3 := DD(13, 34);
		d4 := DD(13, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 41);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 42);
		d2 := DD(13, 43);
		d3 := DD(13, 44);
		d4 := DD(13, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 51);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 52);
		d2 := DD(13, 53);
		d3 := DD(13, 54);
		d4 := DD(13, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 61);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 62);
		d2 := DD(13, 63);
		d3 := DD(13, 64);
		d4 := DD(13, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 71);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 72);
		d2 := DD(13, 73);
		d3 := DD(13, 74);
		d4 := DD(13, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 81);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(13, 82);
		d2 := DD(13, 83);
		d3 := DD(13, 84);
		d4 := DD(13, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(13, 91);
		graph(13, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 12);
		d2 := DD(14, 13);
		d3 := DD(14, 14);
		d4 := DD(14, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 21);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 22);
		d2 := DD(14, 23);
		d3 := DD(14, 24);
		d4 := DD(14, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 31);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 32);
		d2 := DD(14, 33);
		d3 := DD(14, 34);
		d4 := DD(14, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 41);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 42);
		d2 := DD(14, 43);
		d3 := DD(14, 44);
		d4 := DD(14, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 51);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 52);
		d2 := DD(14, 53);
		d3 := DD(14, 54);
		d4 := DD(14, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 61);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 62);
		d2 := DD(14, 63);
		d3 := DD(14, 64);
		d4 := DD(14, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 71);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 72);
		d2 := DD(14, 73);
		d3 := DD(14, 74);
		d4 := DD(14, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 81);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(14, 82);
		d2 := DD(14, 83);
		d3 := DD(14, 84);
		d4 := DD(14, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(14, 91);
		graph(14, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 12);
		d2 := DD(15, 13);
		d3 := DD(15, 14);
		d4 := DD(15, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 21);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 22);
		d2 := DD(15, 23);
		d3 := DD(15, 24);
		d4 := DD(15, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 31);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 32);
		d2 := DD(15, 33);
		d3 := DD(15, 34);
		d4 := DD(15, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 41);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 42);
		d2 := DD(15, 43);
		d3 := DD(15, 44);
		d4 := DD(15, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 51);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 52);
		d2 := DD(15, 53);
		d3 := DD(15, 54);
		d4 := DD(15, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 61);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 62);
		d2 := DD(15, 63);
		d3 := DD(15, 64);
		d4 := DD(15, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 71);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 72);
		d2 := DD(15, 73);
		d3 := DD(15, 74);
		d4 := DD(15, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 81);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(15, 82);
		d2 := DD(15, 83);
		d3 := DD(15, 84);
		d4 := DD(15, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(15, 91);
		graph(15, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 12);
		d2 := DD(16, 13);
		d3 := DD(16, 14);
		d4 := DD(16, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 21);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 22);
		d2 := DD(16, 23);
		d3 := DD(16, 24);
		d4 := DD(16, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 31);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 32);
		d2 := DD(16, 33);
		d3 := DD(16, 34);
		d4 := DD(16, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 41);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 42);
		d2 := DD(16, 43);
		d3 := DD(16, 44);
		d4 := DD(16, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 51);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 52);
		d2 := DD(16, 53);
		d3 := DD(16, 54);
		d4 := DD(16, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 61);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 62);
		d2 := DD(16, 63);
		d3 := DD(16, 64);
		d4 := DD(16, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 71);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 72);
		d2 := DD(16, 73);
		d3 := DD(16, 74);
		d4 := DD(16, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 81);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(16, 82);
		d2 := DD(16, 83);
		d3 := DD(16, 84);
		d4 := DD(16, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(16, 91);
		graph(16, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 12);
		d2 := DD(17, 13);
		d3 := DD(17, 14);
		d4 := DD(17, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 21);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 22);
		d2 := DD(17, 23);
		d3 := DD(17, 24);
		d4 := DD(17, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 31);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 32);
		d2 := DD(17, 33);
		d3 := DD(17, 34);
		d4 := DD(17, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 41);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 42);
		d2 := DD(17, 43);
		d3 := DD(17, 44);
		d4 := DD(17, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 51);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 52);
		d2 := DD(17, 53);
		d3 := DD(17, 54);
		d4 := DD(17, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 61);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 62);
		d2 := DD(17, 63);
		d3 := DD(17, 64);
		d4 := DD(17, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 71);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 72);
		d2 := DD(17, 73);
		d3 := DD(17, 74);
		d4 := DD(17, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 81);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(17, 82);
		d2 := DD(17, 83);
		d3 := DD(17, 84);
		d4 := DD(17, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(17, 91);
		graph(17, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 12);
		d2 := DD(18, 13);
		d3 := DD(18, 14);
		d4 := DD(18, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 21);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 22);
		d2 := DD(18, 23);
		d3 := DD(18, 24);
		d4 := DD(18, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 31);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 32);
		d2 := DD(18, 33);
		d3 := DD(18, 34);
		d4 := DD(18, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 41);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 42);
		d2 := DD(18, 43);
		d3 := DD(18, 44);
		d4 := DD(18, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 51);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 52);
		d2 := DD(18, 53);
		d3 := DD(18, 54);
		d4 := DD(18, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 61);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 62);
		d2 := DD(18, 63);
		d3 := DD(18, 64);
		d4 := DD(18, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 71);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 72);
		d2 := DD(18, 73);
		d3 := DD(18, 74);
		d4 := DD(18, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 81);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(18, 82);
		d2 := DD(18, 83);
		d3 := DD(18, 84);
		d4 := DD(18, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(18, 91);
		graph(18, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 12);
		d2 := DD(19, 13);
		d3 := DD(19, 14);
		d4 := DD(19, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 21);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 22);
		d2 := DD(19, 23);
		d3 := DD(19, 24);
		d4 := DD(19, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 31);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 32);
		d2 := DD(19, 33);
		d3 := DD(19, 34);
		d4 := DD(19, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 41);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 42);
		d2 := DD(19, 43);
		d3 := DD(19, 44);
		d4 := DD(19, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 51);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 52);
		d2 := DD(19, 53);
		d3 := DD(19, 54);
		d4 := DD(19, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 61);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 62);
		d2 := DD(19, 63);
		d3 := DD(19, 64);
		d4 := DD(19, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 71);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 72);
		d2 := DD(19, 73);
		d3 := DD(19, 74);
		d4 := DD(19, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 81);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(19, 82);
		d2 := DD(19, 83);
		d3 := DD(19, 84);
		d4 := DD(19, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(19, 91);
		graph(19, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 12);
		d2 := DD(20, 13);
		d3 := DD(20, 14);
		d4 := DD(20, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 21);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 22);
		d2 := DD(20, 23);
		d3 := DD(20, 24);
		d4 := DD(20, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 31);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 32);
		d2 := DD(20, 33);
		d3 := DD(20, 34);
		d4 := DD(20, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 41);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 42);
		d2 := DD(20, 43);
		d3 := DD(20, 44);
		d4 := DD(20, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 51);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 52);
		d2 := DD(20, 53);
		d3 := DD(20, 54);
		d4 := DD(20, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 61);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 62);
		d2 := DD(20, 63);
		d3 := DD(20, 64);
		d4 := DD(20, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 71);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 72);
		d2 := DD(20, 73);
		d3 := DD(20, 74);
		d4 := DD(20, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 81);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(20, 82);
		d2 := DD(20, 83);
		d3 := DD(20, 84);
		d4 := DD(20, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(20, 91);
		graph(20, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 12);
		d2 := DD(21, 13);
		d3 := DD(21, 14);
		d4 := DD(21, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 21);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 22);
		d2 := DD(21, 23);
		d3 := DD(21, 24);
		d4 := DD(21, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 31);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 32);
		d2 := DD(21, 33);
		d3 := DD(21, 34);
		d4 := DD(21, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 41);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 42);
		d2 := DD(21, 43);
		d3 := DD(21, 44);
		d4 := DD(21, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 51);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 52);
		d2 := DD(21, 53);
		d3 := DD(21, 54);
		d4 := DD(21, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 61);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 62);
		d2 := DD(21, 63);
		d3 := DD(21, 64);
		d4 := DD(21, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 71);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 72);
		d2 := DD(21, 73);
		d3 := DD(21, 74);
		d4 := DD(21, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 81);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(21, 82);
		d2 := DD(21, 83);
		d3 := DD(21, 84);
		d4 := DD(21, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(21, 91);
		graph(21, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 12);
		d2 := DD(22, 13);
		d3 := DD(22, 14);
		d4 := DD(22, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 21);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 22);
		d2 := DD(22, 23);
		d3 := DD(22, 24);
		d4 := DD(22, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 31);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 32);
		d2 := DD(22, 33);
		d3 := DD(22, 34);
		d4 := DD(22, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 41);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 42);
		d2 := DD(22, 43);
		d3 := DD(22, 44);
		d4 := DD(22, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 51);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 52);
		d2 := DD(22, 53);
		d3 := DD(22, 54);
		d4 := DD(22, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 61);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 62);
		d2 := DD(22, 63);
		d3 := DD(22, 64);
		d4 := DD(22, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 71);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 72);
		d2 := DD(22, 73);
		d3 := DD(22, 74);
		d4 := DD(22, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 81);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(22, 82);
		d2 := DD(22, 83);
		d3 := DD(22, 84);
		d4 := DD(22, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(22, 91);
		graph(22, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 12);
		d2 := DD(23, 13);
		d3 := DD(23, 14);
		d4 := DD(23, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 21);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 22);
		d2 := DD(23, 23);
		d3 := DD(23, 24);
		d4 := DD(23, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 31);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 32);
		d2 := DD(23, 33);
		d3 := DD(23, 34);
		d4 := DD(23, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 41);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 42);
		d2 := DD(23, 43);
		d3 := DD(23, 44);
		d4 := DD(23, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 51);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 52);
		d2 := DD(23, 53);
		d3 := DD(23, 54);
		d4 := DD(23, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 61);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 62);
		d2 := DD(23, 63);
		d3 := DD(23, 64);
		d4 := DD(23, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 71);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 72);
		d2 := DD(23, 73);
		d3 := DD(23, 74);
		d4 := DD(23, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 81);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(23, 82);
		d2 := DD(23, 83);
		d3 := DD(23, 84);
		d4 := DD(23, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(23, 91);
		graph(23, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 12);
		d2 := DD(24, 13);
		d3 := DD(24, 14);
		d4 := DD(24, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 21);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 22);
		d2 := DD(24, 23);
		d3 := DD(24, 24);
		d4 := DD(24, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 31);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 32);
		d2 := DD(24, 33);
		d3 := DD(24, 34);
		d4 := DD(24, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 41);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 42);
		d2 := DD(24, 43);
		d3 := DD(24, 44);
		d4 := DD(24, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 51);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 52);
		d2 := DD(24, 53);
		d3 := DD(24, 54);
		d4 := DD(24, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 61);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 62);
		d2 := DD(24, 63);
		d3 := DD(24, 64);
		d4 := DD(24, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 71);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 72);
		d2 := DD(24, 73);
		d3 := DD(24, 74);
		d4 := DD(24, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 81);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(24, 82);
		d2 := DD(24, 83);
		d3 := DD(24, 84);
		d4 := DD(24, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(24, 91);
		graph(24, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 12);
		d2 := DD(25, 13);
		d3 := DD(25, 14);
		d4 := DD(25, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 21);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 22);
		d2 := DD(25, 23);
		d3 := DD(25, 24);
		d4 := DD(25, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 31);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 32);
		d2 := DD(25, 33);
		d3 := DD(25, 34);
		d4 := DD(25, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 41);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 42);
		d2 := DD(25, 43);
		d3 := DD(25, 44);
		d4 := DD(25, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 51);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 52);
		d2 := DD(25, 53);
		d3 := DD(25, 54);
		d4 := DD(25, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 61);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 62);
		d2 := DD(25, 63);
		d3 := DD(25, 64);
		d4 := DD(25, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 71);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 72);
		d2 := DD(25, 73);
		d3 := DD(25, 74);
		d4 := DD(25, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 81);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(25, 82);
		d2 := DD(25, 83);
		d3 := DD(25, 84);
		d4 := DD(25, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(25, 91);
		graph(25, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 12);
		d2 := DD(26, 13);
		d3 := DD(26, 14);
		d4 := DD(26, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 21);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 22);
		d2 := DD(26, 23);
		d3 := DD(26, 24);
		d4 := DD(26, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 31);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 32);
		d2 := DD(26, 33);
		d3 := DD(26, 34);
		d4 := DD(26, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 41);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 42);
		d2 := DD(26, 43);
		d3 := DD(26, 44);
		d4 := DD(26, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 51);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 52);
		d2 := DD(26, 53);
		d3 := DD(26, 54);
		d4 := DD(26, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 61);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 62);
		d2 := DD(26, 63);
		d3 := DD(26, 64);
		d4 := DD(26, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 71);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 72);
		d2 := DD(26, 73);
		d3 := DD(26, 74);
		d4 := DD(26, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 81);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(26, 82);
		d2 := DD(26, 83);
		d3 := DD(26, 84);
		d4 := DD(26, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(26, 91);
		graph(26, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 12);
		d2 := DD(27, 13);
		d3 := DD(27, 14);
		d4 := DD(27, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 21);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 22);
		d2 := DD(27, 23);
		d3 := DD(27, 24);
		d4 := DD(27, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 31);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 32);
		d2 := DD(27, 33);
		d3 := DD(27, 34);
		d4 := DD(27, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 41);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 42);
		d2 := DD(27, 43);
		d3 := DD(27, 44);
		d4 := DD(27, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 51);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 52);
		d2 := DD(27, 53);
		d3 := DD(27, 54);
		d4 := DD(27, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 61);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 62);
		d2 := DD(27, 63);
		d3 := DD(27, 64);
		d4 := DD(27, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 71);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 72);
		d2 := DD(27, 73);
		d3 := DD(27, 74);
		d4 := DD(27, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 81);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(27, 82);
		d2 := DD(27, 83);
		d3 := DD(27, 84);
		d4 := DD(27, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(27, 91);
		graph(27, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 12);
		d2 := DD(28, 13);
		d3 := DD(28, 14);
		d4 := DD(28, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 21);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 22);
		d2 := DD(28, 23);
		d3 := DD(28, 24);
		d4 := DD(28, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 31);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 32);
		d2 := DD(28, 33);
		d3 := DD(28, 34);
		d4 := DD(28, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 41);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 42);
		d2 := DD(28, 43);
		d3 := DD(28, 44);
		d4 := DD(28, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 51);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 52);
		d2 := DD(28, 53);
		d3 := DD(28, 54);
		d4 := DD(28, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 61);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 62);
		d2 := DD(28, 63);
		d3 := DD(28, 64);
		d4 := DD(28, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 71);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 72);
		d2 := DD(28, 73);
		d3 := DD(28, 74);
		d4 := DD(28, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 81);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(28, 82);
		d2 := DD(28, 83);
		d3 := DD(28, 84);
		d4 := DD(28, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(28, 91);
		graph(28, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 12);
		d2 := DD(29, 13);
		d3 := DD(29, 14);
		d4 := DD(29, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 21);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 22);
		d2 := DD(29, 23);
		d3 := DD(29, 24);
		d4 := DD(29, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 31);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 32);
		d2 := DD(29, 33);
		d3 := DD(29, 34);
		d4 := DD(29, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 41);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 42);
		d2 := DD(29, 43);
		d3 := DD(29, 44);
		d4 := DD(29, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 51);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 52);
		d2 := DD(29, 53);
		d3 := DD(29, 54);
		d4 := DD(29, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 61);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 62);
		d2 := DD(29, 63);
		d3 := DD(29, 64);
		d4 := DD(29, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 71);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 72);
		d2 := DD(29, 73);
		d3 := DD(29, 74);
		d4 := DD(29, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 81);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(29, 82);
		d2 := DD(29, 83);
		d3 := DD(29, 84);
		d4 := DD(29, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(29, 91);
		graph(29, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 12);
		d2 := DD(30, 13);
		d3 := DD(30, 14);
		d4 := DD(30, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 21);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 22);
		d2 := DD(30, 23);
		d3 := DD(30, 24);
		d4 := DD(30, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 31);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 32);
		d2 := DD(30, 33);
		d3 := DD(30, 34);
		d4 := DD(30, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 41);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 42);
		d2 := DD(30, 43);
		d3 := DD(30, 44);
		d4 := DD(30, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 51);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 52);
		d2 := DD(30, 53);
		d3 := DD(30, 54);
		d4 := DD(30, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 61);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 62);
		d2 := DD(30, 63);
		d3 := DD(30, 64);
		d4 := DD(30, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 71);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 72);
		d2 := DD(30, 73);
		d3 := DD(30, 74);
		d4 := DD(30, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 81);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(30, 82);
		d2 := DD(30, 83);
		d3 := DD(30, 84);
		d4 := DD(30, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(30, 91);
		graph(30, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 12);
		d2 := DD(31, 13);
		d3 := DD(31, 14);
		d4 := DD(31, 15);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 21);
		graph(31, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 22);
		d2 := DD(31, 23);
		d3 := DD(31, 24);
		d4 := DD(31, 25);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 31);
		graph(31, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 32);
		d2 := DD(31, 33);
		d3 := DD(31, 34);
		d4 := DD(31, 35);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 41);
		graph(31, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 42);
		d2 := DD(31, 43);
		d3 := DD(31, 44);
		d4 := DD(31, 45);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 51);
		graph(31, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 52);
		d2 := DD(31, 53);
		d3 := DD(31, 54);
		d4 := DD(31, 55);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 61);
		graph(31, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 62);
		d2 := DD(31, 63);
		d3 := DD(31, 64);
		d4 := DD(31, 65);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 71);
		graph(31, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 72);
		d2 := DD(31, 73);
		d3 := DD(31, 74);
		d4 := DD(31, 75);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 81);
		graph(31, to_integer(unsigned(d))) <= e2;
		d1 := DD(31, 82);
		d2 := DD(31, 83);
		d3 := DD(31, 84);
		d4 := DD(31, 85);
		d := d1 & d2 & d3 & d4;
		e2 := DD(31, 91);
		graph(31, to_integer(unsigned(d))) <= e2;
		extraction_done <= '1';
	else extraction_done <= '0';
	end if;
	END PROCESS;

END behavioural;