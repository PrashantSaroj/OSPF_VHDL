LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE WORK.ddPackage.ALL;

entity extract_info is
	port(
		DD : in databaseDescription;
		graph: out RAM_FOR_GRAPH:=(others => (others => (others => '1')));
		IP_ADDR : out ip_addr_array);
end extract_info;

architecture behavioural of extract_info is
begin
	-- assumption router ids are 0-31
	IP_ADDR(to_integer(unsigned(DD(0, 4 to 7)))) <= DD(0, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(1, 4 to 7)))) <= DD(1, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(2, 4 to 7)))) <= DD(2, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(3, 4 to 7)))) <= DD(3, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(4, 4 to 7)))) <= DD(4, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(5, 4 to 7)))) <= DD(5, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(6, 4 to 7)))) <= DD(6, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(7, 4 to 7)))) <= DD(7, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(8, 4 to 7)))) <= DD(8, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(9, 4 to 7)))) <= DD(9, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(10, 4 to 7)))) <= DD(10, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(11, 4 to 7)))) <= DD(11, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(12, 4 to 7)))) <= DD(12, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(13, 4 to 7)))) <= DD(13, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(14, 4 to 7)))) <= DD(14, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(15, 4 to 7)))) <= DD(15, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(16, 4 to 7)))) <= DD(16, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(17, 4 to 7)))) <= DD(17, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(18, 4 to 7)))) <= DD(18, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(19, 4 to 7)))) <= DD(19, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(20, 4 to 7)))) <= DD(20, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(21, 4 to 7)))) <= DD(21, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(22, 4 to 7)))) <= DD(22, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(23, 4 to 7)))) <= DD(23, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(24, 4 to 7)))) <= DD(24, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(25, 4 to 7)))) <= DD(25, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(26, 4 to 7)))) <= DD(26, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(27, 4 to 7)))) <= DD(27, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(28, 4 to 7)))) <= DD(28, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(29, 4 to 7)))) <= DD(29, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(30, 4 to 7)))) <= DD(30, 0 to 3);
	IP_ADDR(to_integer(unsigned(DD(31, 4 to 7)))) <= DD(31, 0 to 3);

	-- assigning graph the costs
	graph(0, to_integer(unsigned(DD(0, 12 to 15)))) <= DD(0, 20 to 21);
	graph(0, to_integer(unsigned(DD(0, 22 to 25)))) <= DD(0, 30 to 31);
	graph(0, to_integer(unsigned(DD(0, 32 to 35)))) <= DD(0, 40 to 41);
	graph(0, to_integer(unsigned(DD(0, 42 to 45)))) <= DD(0, 50 to 51);
	graph(0, to_integer(unsigned(DD(0, 52 to 55)))) <= DD(0, 60 to 61);
	graph(0, to_integer(unsigned(DD(0, 62 to 65)))) <= DD(0, 70 to 71);
	graph(0, to_integer(unsigned(DD(0, 72 to 75)))) <= DD(0, 80 to 81);
	graph(0, to_integer(unsigned(DD(0, 82 to 85)))) <= DD(0, 90 to 91);
	graph(1, to_integer(unsigned(DD(1, 12 to 15)))) <= DD(1, 20 to 21);
	graph(1, to_integer(unsigned(DD(1, 22 to 25)))) <= DD(1, 30 to 31);
	graph(1, to_integer(unsigned(DD(1, 32 to 35)))) <= DD(1, 40 to 41);
	graph(1, to_integer(unsigned(DD(1, 42 to 45)))) <= DD(1, 50 to 51);
	graph(1, to_integer(unsigned(DD(1, 52 to 55)))) <= DD(1, 60 to 61);
	graph(1, to_integer(unsigned(DD(1, 62 to 65)))) <= DD(1, 70 to 71);
	graph(1, to_integer(unsigned(DD(1, 72 to 75)))) <= DD(1, 80 to 81);
	graph(1, to_integer(unsigned(DD(1, 82 to 85)))) <= DD(1, 90 to 91);
	graph(2, to_integer(unsigned(DD(2, 12 to 15)))) <= DD(2, 20 to 21);
	graph(2, to_integer(unsigned(DD(2, 22 to 25)))) <= DD(2, 30 to 31);
	graph(2, to_integer(unsigned(DD(2, 32 to 35)))) <= DD(2, 40 to 41);
	graph(2, to_integer(unsigned(DD(2, 42 to 45)))) <= DD(2, 50 to 51);
	graph(2, to_integer(unsigned(DD(2, 52 to 55)))) <= DD(2, 60 to 61);
	graph(2, to_integer(unsigned(DD(2, 62 to 65)))) <= DD(2, 70 to 71);
	graph(2, to_integer(unsigned(DD(2, 72 to 75)))) <= DD(2, 80 to 81);
	graph(2, to_integer(unsigned(DD(2, 82 to 85)))) <= DD(2, 90 to 91);
	graph(3, to_integer(unsigned(DD(3, 12 to 15)))) <= DD(3, 20 to 21);
	graph(3, to_integer(unsigned(DD(3, 22 to 25)))) <= DD(3, 30 to 31);
	graph(3, to_integer(unsigned(DD(3, 32 to 35)))) <= DD(3, 40 to 41);
	graph(3, to_integer(unsigned(DD(3, 42 to 45)))) <= DD(3, 50 to 51);
	graph(3, to_integer(unsigned(DD(3, 52 to 55)))) <= DD(3, 60 to 61);
	graph(3, to_integer(unsigned(DD(3, 62 to 65)))) <= DD(3, 70 to 71);
	graph(3, to_integer(unsigned(DD(3, 72 to 75)))) <= DD(3, 80 to 81);
	graph(3, to_integer(unsigned(DD(3, 82 to 85)))) <= DD(3, 90 to 91);
	graph(4, to_integer(unsigned(DD(4, 12 to 15)))) <= DD(4, 20 to 21);
	graph(4, to_integer(unsigned(DD(4, 22 to 25)))) <= DD(4, 30 to 31);
	graph(4, to_integer(unsigned(DD(4, 32 to 35)))) <= DD(4, 40 to 41);
	graph(4, to_integer(unsigned(DD(4, 42 to 45)))) <= DD(4, 50 to 51);
	graph(4, to_integer(unsigned(DD(4, 52 to 55)))) <= DD(4, 60 to 61);
	graph(4, to_integer(unsigned(DD(4, 62 to 65)))) <= DD(4, 70 to 71);
	graph(4, to_integer(unsigned(DD(4, 72 to 75)))) <= DD(4, 80 to 81);
	graph(4, to_integer(unsigned(DD(4, 82 to 85)))) <= DD(4, 90 to 91);
	graph(5, to_integer(unsigned(DD(5, 12 to 15)))) <= DD(5, 20 to 21);
	graph(5, to_integer(unsigned(DD(5, 22 to 25)))) <= DD(5, 30 to 31);
	graph(5, to_integer(unsigned(DD(5, 32 to 35)))) <= DD(5, 40 to 41);
	graph(5, to_integer(unsigned(DD(5, 42 to 45)))) <= DD(5, 50 to 51);
	graph(5, to_integer(unsigned(DD(5, 52 to 55)))) <= DD(5, 60 to 61);
	graph(5, to_integer(unsigned(DD(5, 62 to 65)))) <= DD(5, 70 to 71);
	graph(5, to_integer(unsigned(DD(5, 72 to 75)))) <= DD(5, 80 to 81);
	graph(5, to_integer(unsigned(DD(5, 82 to 85)))) <= DD(5, 90 to 91);
	graph(6, to_integer(unsigned(DD(6, 12 to 15)))) <= DD(6, 20 to 21);
	graph(6, to_integer(unsigned(DD(6, 22 to 25)))) <= DD(6, 30 to 31);
	graph(6, to_integer(unsigned(DD(6, 32 to 35)))) <= DD(6, 40 to 41);
	graph(6, to_integer(unsigned(DD(6, 42 to 45)))) <= DD(6, 50 to 51);
	graph(6, to_integer(unsigned(DD(6, 52 to 55)))) <= DD(6, 60 to 61);
	graph(6, to_integer(unsigned(DD(6, 62 to 65)))) <= DD(6, 70 to 71);
	graph(6, to_integer(unsigned(DD(6, 72 to 75)))) <= DD(6, 80 to 81);
	graph(6, to_integer(unsigned(DD(6, 82 to 85)))) <= DD(6, 90 to 91);
	graph(7, to_integer(unsigned(DD(7, 12 to 15)))) <= DD(7, 20 to 21);
	graph(7, to_integer(unsigned(DD(7, 22 to 25)))) <= DD(7, 30 to 31);
	graph(7, to_integer(unsigned(DD(7, 32 to 35)))) <= DD(7, 40 to 41);
	graph(7, to_integer(unsigned(DD(7, 42 to 45)))) <= DD(7, 50 to 51);
	graph(7, to_integer(unsigned(DD(7, 52 to 55)))) <= DD(7, 60 to 61);
	graph(7, to_integer(unsigned(DD(7, 62 to 65)))) <= DD(7, 70 to 71);
	graph(7, to_integer(unsigned(DD(7, 72 to 75)))) <= DD(7, 80 to 81);
	graph(7, to_integer(unsigned(DD(7, 82 to 85)))) <= DD(7, 90 to 91);
	graph(8, to_integer(unsigned(DD(8, 12 to 15)))) <= DD(8, 20 to 21);
	graph(8, to_integer(unsigned(DD(8, 22 to 25)))) <= DD(8, 30 to 31);
	graph(8, to_integer(unsigned(DD(8, 32 to 35)))) <= DD(8, 40 to 41);
	graph(8, to_integer(unsigned(DD(8, 42 to 45)))) <= DD(8, 50 to 51);
	graph(8, to_integer(unsigned(DD(8, 52 to 55)))) <= DD(8, 60 to 61);
	graph(8, to_integer(unsigned(DD(8, 62 to 65)))) <= DD(8, 70 to 71);
	graph(8, to_integer(unsigned(DD(8, 72 to 75)))) <= DD(8, 80 to 81);
	graph(8, to_integer(unsigned(DD(8, 82 to 85)))) <= DD(8, 90 to 91);
	graph(9, to_integer(unsigned(DD(9, 12 to 15)))) <= DD(9, 20 to 21);
	graph(9, to_integer(unsigned(DD(9, 22 to 25)))) <= DD(9, 30 to 31);
	graph(9, to_integer(unsigned(DD(9, 32 to 35)))) <= DD(9, 40 to 41);
	graph(9, to_integer(unsigned(DD(9, 42 to 45)))) <= DD(9, 50 to 51);
	graph(9, to_integer(unsigned(DD(9, 52 to 55)))) <= DD(9, 60 to 61);
	graph(9, to_integer(unsigned(DD(9, 62 to 65)))) <= DD(9, 70 to 71);
	graph(9, to_integer(unsigned(DD(9, 72 to 75)))) <= DD(9, 80 to 81);
	graph(9, to_integer(unsigned(DD(9, 82 to 85)))) <= DD(9, 90 to 91);
	graph(10, to_integer(unsigned(DD(10, 12 to 15)))) <= DD(10, 20 to 21);
	graph(10, to_integer(unsigned(DD(10, 22 to 25)))) <= DD(10, 30 to 31);
	graph(10, to_integer(unsigned(DD(10, 32 to 35)))) <= DD(10, 40 to 41);
	graph(10, to_integer(unsigned(DD(10, 42 to 45)))) <= DD(10, 50 to 51);
	graph(10, to_integer(unsigned(DD(10, 52 to 55)))) <= DD(10, 60 to 61);
	graph(10, to_integer(unsigned(DD(10, 62 to 65)))) <= DD(10, 70 to 71);
	graph(10, to_integer(unsigned(DD(10, 72 to 75)))) <= DD(10, 80 to 81);
	graph(10, to_integer(unsigned(DD(10, 82 to 85)))) <= DD(10, 90 to 91);
	graph(11, to_integer(unsigned(DD(11, 12 to 15)))) <= DD(11, 20 to 21);
	graph(11, to_integer(unsigned(DD(11, 22 to 25)))) <= DD(11, 30 to 31);
	graph(11, to_integer(unsigned(DD(11, 32 to 35)))) <= DD(11, 40 to 41);
	graph(11, to_integer(unsigned(DD(11, 42 to 45)))) <= DD(11, 50 to 51);
	graph(11, to_integer(unsigned(DD(11, 52 to 55)))) <= DD(11, 60 to 61);
	graph(11, to_integer(unsigned(DD(11, 62 to 65)))) <= DD(11, 70 to 71);
	graph(11, to_integer(unsigned(DD(11, 72 to 75)))) <= DD(11, 80 to 81);
	graph(11, to_integer(unsigned(DD(11, 82 to 85)))) <= DD(11, 90 to 91);
	graph(12, to_integer(unsigned(DD(12, 12 to 15)))) <= DD(12, 20 to 21);
	graph(12, to_integer(unsigned(DD(12, 22 to 25)))) <= DD(12, 30 to 31);
	graph(12, to_integer(unsigned(DD(12, 32 to 35)))) <= DD(12, 40 to 41);
	graph(12, to_integer(unsigned(DD(12, 42 to 45)))) <= DD(12, 50 to 51);
	graph(12, to_integer(unsigned(DD(12, 52 to 55)))) <= DD(12, 60 to 61);
	graph(12, to_integer(unsigned(DD(12, 62 to 65)))) <= DD(12, 70 to 71);
	graph(12, to_integer(unsigned(DD(12, 72 to 75)))) <= DD(12, 80 to 81);
	graph(12, to_integer(unsigned(DD(12, 82 to 85)))) <= DD(12, 90 to 91);
	graph(13, to_integer(unsigned(DD(13, 12 to 15)))) <= DD(13, 20 to 21);
	graph(13, to_integer(unsigned(DD(13, 22 to 25)))) <= DD(13, 30 to 31);
	graph(13, to_integer(unsigned(DD(13, 32 to 35)))) <= DD(13, 40 to 41);
	graph(13, to_integer(unsigned(DD(13, 42 to 45)))) <= DD(13, 50 to 51);
	graph(13, to_integer(unsigned(DD(13, 52 to 55)))) <= DD(13, 60 to 61);
	graph(13, to_integer(unsigned(DD(13, 62 to 65)))) <= DD(13, 70 to 71);
	graph(13, to_integer(unsigned(DD(13, 72 to 75)))) <= DD(13, 80 to 81);
	graph(13, to_integer(unsigned(DD(13, 82 to 85)))) <= DD(13, 90 to 91);
	graph(14, to_integer(unsigned(DD(14, 12 to 15)))) <= DD(14, 20 to 21);
	graph(14, to_integer(unsigned(DD(14, 22 to 25)))) <= DD(14, 30 to 31);
	graph(14, to_integer(unsigned(DD(14, 32 to 35)))) <= DD(14, 40 to 41);
	graph(14, to_integer(unsigned(DD(14, 42 to 45)))) <= DD(14, 50 to 51);
	graph(14, to_integer(unsigned(DD(14, 52 to 55)))) <= DD(14, 60 to 61);
	graph(14, to_integer(unsigned(DD(14, 62 to 65)))) <= DD(14, 70 to 71);
	graph(14, to_integer(unsigned(DD(14, 72 to 75)))) <= DD(14, 80 to 81);
	graph(14, to_integer(unsigned(DD(14, 82 to 85)))) <= DD(14, 90 to 91);
	graph(15, to_integer(unsigned(DD(15, 12 to 15)))) <= DD(15, 20 to 21);
	graph(15, to_integer(unsigned(DD(15, 22 to 25)))) <= DD(15, 30 to 31);
	graph(15, to_integer(unsigned(DD(15, 32 to 35)))) <= DD(15, 40 to 41);
	graph(15, to_integer(unsigned(DD(15, 42 to 45)))) <= DD(15, 50 to 51);
	graph(15, to_integer(unsigned(DD(15, 52 to 55)))) <= DD(15, 60 to 61);
	graph(15, to_integer(unsigned(DD(15, 62 to 65)))) <= DD(15, 70 to 71);
	graph(15, to_integer(unsigned(DD(15, 72 to 75)))) <= DD(15, 80 to 81);
	graph(15, to_integer(unsigned(DD(15, 82 to 85)))) <= DD(15, 90 to 91);
	graph(16, to_integer(unsigned(DD(16, 12 to 15)))) <= DD(16, 20 to 21);
	graph(16, to_integer(unsigned(DD(16, 22 to 25)))) <= DD(16, 30 to 31);
	graph(16, to_integer(unsigned(DD(16, 32 to 35)))) <= DD(16, 40 to 41);
	graph(16, to_integer(unsigned(DD(16, 42 to 45)))) <= DD(16, 50 to 51);
	graph(16, to_integer(unsigned(DD(16, 52 to 55)))) <= DD(16, 60 to 61);
	graph(16, to_integer(unsigned(DD(16, 62 to 65)))) <= DD(16, 70 to 71);
	graph(16, to_integer(unsigned(DD(16, 72 to 75)))) <= DD(16, 80 to 81);
	graph(16, to_integer(unsigned(DD(16, 82 to 85)))) <= DD(16, 90 to 91);
	graph(17, to_integer(unsigned(DD(17, 12 to 15)))) <= DD(17, 20 to 21);
	graph(17, to_integer(unsigned(DD(17, 22 to 25)))) <= DD(17, 30 to 31);
	graph(17, to_integer(unsigned(DD(17, 32 to 35)))) <= DD(17, 40 to 41);
	graph(17, to_integer(unsigned(DD(17, 42 to 45)))) <= DD(17, 50 to 51);
	graph(17, to_integer(unsigned(DD(17, 52 to 55)))) <= DD(17, 60 to 61);
	graph(17, to_integer(unsigned(DD(17, 62 to 65)))) <= DD(17, 70 to 71);
	graph(17, to_integer(unsigned(DD(17, 72 to 75)))) <= DD(17, 80 to 81);
	graph(17, to_integer(unsigned(DD(17, 82 to 85)))) <= DD(17, 90 to 91);
	graph(18, to_integer(unsigned(DD(18, 12 to 15)))) <= DD(18, 20 to 21);
	graph(18, to_integer(unsigned(DD(18, 22 to 25)))) <= DD(18, 30 to 31);
	graph(18, to_integer(unsigned(DD(18, 32 to 35)))) <= DD(18, 40 to 41);
	graph(18, to_integer(unsigned(DD(18, 42 to 45)))) <= DD(18, 50 to 51);
	graph(18, to_integer(unsigned(DD(18, 52 to 55)))) <= DD(18, 60 to 61);
	graph(18, to_integer(unsigned(DD(18, 62 to 65)))) <= DD(18, 70 to 71);
	graph(18, to_integer(unsigned(DD(18, 72 to 75)))) <= DD(18, 80 to 81);
	graph(18, to_integer(unsigned(DD(18, 82 to 85)))) <= DD(18, 90 to 91);
	graph(19, to_integer(unsigned(DD(19, 12 to 15)))) <= DD(19, 20 to 21);
	graph(19, to_integer(unsigned(DD(19, 22 to 25)))) <= DD(19, 30 to 31);
	graph(19, to_integer(unsigned(DD(19, 32 to 35)))) <= DD(19, 40 to 41);
	graph(19, to_integer(unsigned(DD(19, 42 to 45)))) <= DD(19, 50 to 51);
	graph(19, to_integer(unsigned(DD(19, 52 to 55)))) <= DD(19, 60 to 61);
	graph(19, to_integer(unsigned(DD(19, 62 to 65)))) <= DD(19, 70 to 71);
	graph(19, to_integer(unsigned(DD(19, 72 to 75)))) <= DD(19, 80 to 81);
	graph(19, to_integer(unsigned(DD(19, 82 to 85)))) <= DD(19, 90 to 91);
	graph(20, to_integer(unsigned(DD(20, 12 to 15)))) <= DD(20, 20 to 21);
	graph(20, to_integer(unsigned(DD(20, 22 to 25)))) <= DD(20, 30 to 31);
	graph(20, to_integer(unsigned(DD(20, 32 to 35)))) <= DD(20, 40 to 41);
	graph(20, to_integer(unsigned(DD(20, 42 to 45)))) <= DD(20, 50 to 51);
	graph(20, to_integer(unsigned(DD(20, 52 to 55)))) <= DD(20, 60 to 61);
	graph(20, to_integer(unsigned(DD(20, 62 to 65)))) <= DD(20, 70 to 71);
	graph(20, to_integer(unsigned(DD(20, 72 to 75)))) <= DD(20, 80 to 81);
	graph(20, to_integer(unsigned(DD(20, 82 to 85)))) <= DD(20, 90 to 91);
	graph(21, to_integer(unsigned(DD(21, 12 to 15)))) <= DD(21, 20 to 21);
	graph(21, to_integer(unsigned(DD(21, 22 to 25)))) <= DD(21, 30 to 31);
	graph(21, to_integer(unsigned(DD(21, 32 to 35)))) <= DD(21, 40 to 41);
	graph(21, to_integer(unsigned(DD(21, 42 to 45)))) <= DD(21, 50 to 51);
	graph(21, to_integer(unsigned(DD(21, 52 to 55)))) <= DD(21, 60 to 61);
	graph(21, to_integer(unsigned(DD(21, 62 to 65)))) <= DD(21, 70 to 71);
	graph(21, to_integer(unsigned(DD(21, 72 to 75)))) <= DD(21, 80 to 81);
	graph(21, to_integer(unsigned(DD(21, 82 to 85)))) <= DD(21, 90 to 91);
	graph(22, to_integer(unsigned(DD(22, 12 to 15)))) <= DD(22, 20 to 21);
	graph(22, to_integer(unsigned(DD(22, 22 to 25)))) <= DD(22, 30 to 31);
	graph(22, to_integer(unsigned(DD(22, 32 to 35)))) <= DD(22, 40 to 41);
	graph(22, to_integer(unsigned(DD(22, 42 to 45)))) <= DD(22, 50 to 51);
	graph(22, to_integer(unsigned(DD(22, 52 to 55)))) <= DD(22, 60 to 61);
	graph(22, to_integer(unsigned(DD(22, 62 to 65)))) <= DD(22, 70 to 71);
	graph(22, to_integer(unsigned(DD(22, 72 to 75)))) <= DD(22, 80 to 81);
	graph(22, to_integer(unsigned(DD(22, 82 to 85)))) <= DD(22, 90 to 91);
	graph(23, to_integer(unsigned(DD(23, 12 to 15)))) <= DD(23, 20 to 21);
	graph(23, to_integer(unsigned(DD(23, 22 to 25)))) <= DD(23, 30 to 31);
	graph(23, to_integer(unsigned(DD(23, 32 to 35)))) <= DD(23, 40 to 41);
	graph(23, to_integer(unsigned(DD(23, 42 to 45)))) <= DD(23, 50 to 51);
	graph(23, to_integer(unsigned(DD(23, 52 to 55)))) <= DD(23, 60 to 61);
	graph(23, to_integer(unsigned(DD(23, 62 to 65)))) <= DD(23, 70 to 71);
	graph(23, to_integer(unsigned(DD(23, 72 to 75)))) <= DD(23, 80 to 81);
	graph(23, to_integer(unsigned(DD(23, 82 to 85)))) <= DD(23, 90 to 91);
	graph(24, to_integer(unsigned(DD(24, 12 to 15)))) <= DD(24, 20 to 21);
	graph(24, to_integer(unsigned(DD(24, 22 to 25)))) <= DD(24, 30 to 31);
	graph(24, to_integer(unsigned(DD(24, 32 to 35)))) <= DD(24, 40 to 41);
	graph(24, to_integer(unsigned(DD(24, 42 to 45)))) <= DD(24, 50 to 51);
	graph(24, to_integer(unsigned(DD(24, 52 to 55)))) <= DD(24, 60 to 61);
	graph(24, to_integer(unsigned(DD(24, 62 to 65)))) <= DD(24, 70 to 71);
	graph(24, to_integer(unsigned(DD(24, 72 to 75)))) <= DD(24, 80 to 81);
	graph(24, to_integer(unsigned(DD(24, 82 to 85)))) <= DD(24, 90 to 91);
	graph(25, to_integer(unsigned(DD(25, 12 to 15)))) <= DD(25, 20 to 21);
	graph(25, to_integer(unsigned(DD(25, 22 to 25)))) <= DD(25, 30 to 31);
	graph(25, to_integer(unsigned(DD(25, 32 to 35)))) <= DD(25, 40 to 41);
	graph(25, to_integer(unsigned(DD(25, 42 to 45)))) <= DD(25, 50 to 51);
	graph(25, to_integer(unsigned(DD(25, 52 to 55)))) <= DD(25, 60 to 61);
	graph(25, to_integer(unsigned(DD(25, 62 to 65)))) <= DD(25, 70 to 71);
	graph(25, to_integer(unsigned(DD(25, 72 to 75)))) <= DD(25, 80 to 81);
	graph(25, to_integer(unsigned(DD(25, 82 to 85)))) <= DD(25, 90 to 91);
	graph(26, to_integer(unsigned(DD(26, 12 to 15)))) <= DD(26, 20 to 21);
	graph(26, to_integer(unsigned(DD(26, 22 to 25)))) <= DD(26, 30 to 31);
	graph(26, to_integer(unsigned(DD(26, 32 to 35)))) <= DD(26, 40 to 41);
	graph(26, to_integer(unsigned(DD(26, 42 to 45)))) <= DD(26, 50 to 51);
	graph(26, to_integer(unsigned(DD(26, 52 to 55)))) <= DD(26, 60 to 61);
	graph(26, to_integer(unsigned(DD(26, 62 to 65)))) <= DD(26, 70 to 71);
	graph(26, to_integer(unsigned(DD(26, 72 to 75)))) <= DD(26, 80 to 81);
	graph(26, to_integer(unsigned(DD(26, 82 to 85)))) <= DD(26, 90 to 91);
	graph(27, to_integer(unsigned(DD(27, 12 to 15)))) <= DD(27, 20 to 21);
	graph(27, to_integer(unsigned(DD(27, 22 to 25)))) <= DD(27, 30 to 31);
	graph(27, to_integer(unsigned(DD(27, 32 to 35)))) <= DD(27, 40 to 41);
	graph(27, to_integer(unsigned(DD(27, 42 to 45)))) <= DD(27, 50 to 51);
	graph(27, to_integer(unsigned(DD(27, 52 to 55)))) <= DD(27, 60 to 61);
	graph(27, to_integer(unsigned(DD(27, 62 to 65)))) <= DD(27, 70 to 71);
	graph(27, to_integer(unsigned(DD(27, 72 to 75)))) <= DD(27, 80 to 81);
	graph(27, to_integer(unsigned(DD(27, 82 to 85)))) <= DD(27, 90 to 91);
	graph(28, to_integer(unsigned(DD(28, 12 to 15)))) <= DD(28, 20 to 21);
	graph(28, to_integer(unsigned(DD(28, 22 to 25)))) <= DD(28, 30 to 31);
	graph(28, to_integer(unsigned(DD(28, 32 to 35)))) <= DD(28, 40 to 41);
	graph(28, to_integer(unsigned(DD(28, 42 to 45)))) <= DD(28, 50 to 51);
	graph(28, to_integer(unsigned(DD(28, 52 to 55)))) <= DD(28, 60 to 61);
	graph(28, to_integer(unsigned(DD(28, 62 to 65)))) <= DD(28, 70 to 71);
	graph(28, to_integer(unsigned(DD(28, 72 to 75)))) <= DD(28, 80 to 81);
	graph(28, to_integer(unsigned(DD(28, 82 to 85)))) <= DD(28, 90 to 91);
	graph(29, to_integer(unsigned(DD(29, 12 to 15)))) <= DD(29, 20 to 21);
	graph(29, to_integer(unsigned(DD(29, 22 to 25)))) <= DD(29, 30 to 31);
	graph(29, to_integer(unsigned(DD(29, 32 to 35)))) <= DD(29, 40 to 41);
	graph(29, to_integer(unsigned(DD(29, 42 to 45)))) <= DD(29, 50 to 51);
	graph(29, to_integer(unsigned(DD(29, 52 to 55)))) <= DD(29, 60 to 61);
	graph(29, to_integer(unsigned(DD(29, 62 to 65)))) <= DD(29, 70 to 71);
	graph(29, to_integer(unsigned(DD(29, 72 to 75)))) <= DD(29, 80 to 81);
	graph(29, to_integer(unsigned(DD(29, 82 to 85)))) <= DD(29, 90 to 91);
	graph(30, to_integer(unsigned(DD(30, 12 to 15)))) <= DD(30, 20 to 21);
	graph(30, to_integer(unsigned(DD(30, 22 to 25)))) <= DD(30, 30 to 31);
	graph(30, to_integer(unsigned(DD(30, 32 to 35)))) <= DD(30, 40 to 41);
	graph(30, to_integer(unsigned(DD(30, 42 to 45)))) <= DD(30, 50 to 51);
	graph(30, to_integer(unsigned(DD(30, 52 to 55)))) <= DD(30, 60 to 61);
	graph(30, to_integer(unsigned(DD(30, 62 to 65)))) <= DD(30, 70 to 71);
	graph(30, to_integer(unsigned(DD(30, 72 to 75)))) <= DD(30, 80 to 81);
	graph(30, to_integer(unsigned(DD(30, 82 to 85)))) <= DD(30, 90 to 91);
	graph(31, to_integer(unsigned(DD(31, 12 to 15)))) <= DD(31, 20 to 21);
	graph(31, to_integer(unsigned(DD(31, 22 to 25)))) <= DD(31, 30 to 31);
	graph(31, to_integer(unsigned(DD(31, 32 to 35)))) <= DD(31, 40 to 41);
	graph(31, to_integer(unsigned(DD(31, 42 to 45)))) <= DD(31, 50 to 51);
	graph(31, to_integer(unsigned(DD(31, 52 to 55)))) <= DD(31, 60 to 61);
	graph(31, to_integer(unsigned(DD(31, 62 to 65)))) <= DD(31, 70 to 71);
	graph(31, to_integer(unsigned(DD(31, 72 to 75)))) <= DD(31, 80 to 81);
	graph(31, to_integer(unsigned(DD(31, 82 to 85)))) <= DD(31, 90 to 91);
end behavioural;
