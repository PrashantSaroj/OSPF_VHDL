-- TestBench Template 
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY tb_dd IS
END tb_dd;
ARCHITECTURE behavior OF tb_dd IS 
-- Component Declaration
        COMPONENT ans_lsReq
        PORT(
                clk: in std_logic;
                packet_in1: in std_logic_vector(7 downto 0);
                valid_in1: in std_logic;
                op: out std_logic_vector(7 downto 0):= "000000000";
                is_op: out std_logic:= '0';
                graph: in RAM_FOR_GRAPH
                );
        END COMPONENT;
          
          signal clk: std_logic := '0';
        SIGNAL packet_in1 :  std_logic_vector(7 downto 0);
        SIGNAL valid_in1 : std_logic;

        signal op: std_logic_vector(7 downto 0):= "000000000";
        signal graph: RAM_FOR_GRAPH;
        signal is_op: std_logic:= '0';
        
           -- Clock period definitions
 constant clk_period : time := 10 ns;
BEGIN
      
-- Component Instantiation
        uut: ans_lsReq PORT MAP(
                clk => clk,
                packet_in => packet_in1,
                valid_in => valid_in1,
                op => op,
                graph => graph,
                is_op => is_op
        );

        clk_process :process
begin
clk <= '0';
wait for clk_period/2;
clk <= '1';
wait for clk_period/2;
end process;

--  Test Bench Statements
   tb : PROCESS
   BEGIN
    -- wait until global set/reset completes
    -- Add user defined stimulus here
    valid_in1 <= '1';

    graph(0,0) <= "11111111"
    graph(0,1) <= "11111111"
    graph(0,2) <= "11111111"
    graph(0,3) <= "11111111"
    graph(0,4) <= "11111111"
    graph(0,5) <= "11111111"
    graph(0,6) <= "11111111"
    graph(0,7) <= "11111111"
    graph(0,8) <= "11111111"
    graph(0,9) <= "11111111"
    graph(0,10) <= "11111111"
    graph(0,11) <= "11111111"
    graph(0,12) <= "11111111"
    graph(0,13) <= "11111111"
    graph(0,14) <= "11111111"
    graph(0,15) <= "11111111"
    graph(0,16) <= "11111111"
    graph(0,17) <= "11111111"
    graph(0,18) <= "11111111"
    graph(0,19) <= "11111111"
    graph(0,20) <= "11111111"
    graph(0,21) <= "11111111"
    graph(0,22) <= "11111111"
    graph(0,23) <= "11111111"
    graph(0,24) <= "11111111"
    graph(0,25) <= "11111111"
    graph(0,26) <= "11111111"
    graph(0,27) <= "11111111"
    graph(0,28) <= "11111111"
    graph(0,29) <= "11111111"
    graph(0,30) <= "11111111"
    graph(0,31) <= "11111111"
    graph(1,0) <= "11111111"
    graph(1,1) <= "11111111"
    graph(1,2) <= "11111111"
    graph(1,3) <= "11111111"
    graph(1,4) <= "11111111"
    graph(1,5) <= "11111111"
    graph(1,6) <= "11111111"
    graph(1,7) <= "11111111"
    graph(1,8) <= "11111111"
    graph(1,9) <= "11111111"
    graph(1,10) <= "11111111"
    graph(1,11) <= "11111111"
    graph(1,12) <= "11111111"
    graph(1,13) <= "11111111"
    graph(1,14) <= "11111111"
    graph(1,15) <= "11111111"
    graph(1,16) <= "11111111"
    graph(1,17) <= "11111111"
    graph(1,18) <= "11111111"
    graph(1,19) <= "11111111"
    graph(1,20) <= "11111111"
    graph(1,21) <= "11111111"
    graph(1,22) <= "11111111"
    graph(1,23) <= "11111111"
    graph(1,24) <= "11111111"
    graph(1,25) <= "11111111"
    graph(1,26) <= "11111111"
    graph(1,27) <= "11111111"
    graph(1,28) <= "11111111"
    graph(1,29) <= "11111111"
    graph(1,30) <= "11111111"
    graph(1,31) <= "11111111"
    graph(2,0) <= "11111111"
    graph(2,1) <= "11111111"
    graph(2,2) <= "11111111"
    graph(2,3) <= "11111111"
    graph(2,4) <= "11111111"
    graph(2,5) <= "11111111"
    graph(2,6) <= "11111111"
    graph(2,7) <= "11111111"
    graph(2,8) <= "11111111"
    graph(2,9) <= "11111111"
    graph(2,10) <= "11111111"
    graph(2,11) <= "11111111"
    graph(2,12) <= "11111111"
    graph(2,13) <= "11111111"
    graph(2,14) <= "11111111"
    graph(2,15) <= "11111111"
    graph(2,16) <= "11111111"
    graph(2,17) <= "11111111"
    graph(2,18) <= "11111111"
    graph(2,19) <= "11111111"
    graph(2,20) <= "11111111"
    graph(2,21) <= "11111111"
    graph(2,22) <= "11111111"
    graph(2,23) <= "11111111"
    graph(2,24) <= "11111111"
    graph(2,25) <= "11111111"
    graph(2,26) <= "11111111"
    graph(2,27) <= "11111111"
    graph(2,28) <= "11111111"
    graph(2,29) <= "11111111"
    graph(2,30) <= "11111111"
    graph(2,31) <= "11111111"
    graph(3,0) <= "11111111"
    graph(3,1) <= "11111111"
    graph(3,2) <= "11111111"
    graph(3,3) <= "11111111"
    graph(3,4) <= "11111111"
    graph(3,5) <= "11111111"
    graph(3,6) <= "11111111"
    graph(3,7) <= "11111111"
    graph(3,8) <= "11111111"
    graph(3,9) <= "11111111"
    graph(3,10) <= "11111111"
    graph(3,11) <= "11111111"
    graph(3,12) <= "11111111"
    graph(3,13) <= "11111111"
    graph(3,14) <= "11111111"
    graph(3,15) <= "11111111"
    graph(3,16) <= "11111111"
    graph(3,17) <= "11111111"
    graph(3,18) <= "11111111"
    graph(3,19) <= "11111111"
    graph(3,20) <= "11111111"
    graph(3,21) <= "11111111"
    graph(3,22) <= "11111111"
    graph(3,23) <= "11111111"
    graph(3,24) <= "11111111"
    graph(3,25) <= "11111111"
    graph(3,26) <= "11111111"
    graph(3,27) <= "11111111"
    graph(3,28) <= "11111111"
    graph(3,29) <= "11111111"
    graph(3,30) <= "11111111"
    graph(3,31) <= "11111111"
    graph(4,0) <= "11111111"
    graph(4,1) <= "11111111"
    graph(4,2) <= "11111111"
    graph(4,3) <= "11111111"
    graph(4,4) <= "11111111"
    graph(4,5) <= "11111111"
    graph(4,6) <= "11111111"
    graph(4,7) <= "11111111"
    graph(4,8) <= "11111111"
    graph(4,9) <= "11111111"
    graph(4,10) <= "11111111"
    graph(4,11) <= "11111111"
    graph(4,12) <= "11111111"
    graph(4,13) <= "11111111"
    graph(4,14) <= "11111111"
    graph(4,15) <= "11111111"
    graph(4,16) <= "11111111"
    graph(4,17) <= "11111111"
    graph(4,18) <= "11111111"
    graph(4,19) <= "11111111"
    graph(4,20) <= "11111111"
    graph(4,21) <= "11111111"
    graph(4,22) <= "11111111"
    graph(4,23) <= "11111111"
    graph(4,24) <= "11111111"
    graph(4,25) <= "11111111"
    graph(4,26) <= "11111111"
    graph(4,27) <= "11111111"
    graph(4,28) <= "11111111"
    graph(4,29) <= "11111111"
    graph(4,30) <= "11111111"
    graph(4,31) <= "11111111"
    graph(5,0) <= "11111111"
    graph(5,1) <= "11111111"
    graph(5,2) <= "11111111"
    graph(5,3) <= "11111111"
    graph(5,4) <= "11111111"
    graph(5,5) <= "11111111"
    graph(5,6) <= "11111111"
    graph(5,7) <= "11111111"
    graph(5,8) <= "11111111"
    graph(5,9) <= "11111111"
    graph(5,10) <= "11111111"
    graph(5,11) <= "11111111"
    graph(5,12) <= "11111111"
    graph(5,13) <= "11111111"
    graph(5,14) <= "11111111"
    graph(5,15) <= "11111111"
    graph(5,16) <= "11111111"
    graph(5,17) <= "11111111"
    graph(5,18) <= "11111111"
    graph(5,19) <= "11111111"
    graph(5,20) <= "11111111"
    graph(5,21) <= "11111111"
    graph(5,22) <= "11111111"
    graph(5,23) <= "11111111"
    graph(5,24) <= "11111111"
    graph(5,25) <= "11111111"
    graph(5,26) <= "11111111"
    graph(5,27) <= "11111111"
    graph(5,28) <= "11111111"
    graph(5,29) <= "11111111"
    graph(5,30) <= "11111111"
    graph(5,31) <= "11111111"
    graph(6,0) <= "11111111"
    graph(6,1) <= "11111111"
    graph(6,2) <= "11111111"
    graph(6,3) <= "11111111"
    graph(6,4) <= "11111111"
    graph(6,5) <= "11111111"
    graph(6,6) <= "11111111"
    graph(6,7) <= "11111111"
    graph(6,8) <= "11111111"
    graph(6,9) <= "11111111"
    graph(6,10) <= "11111111"
    graph(6,11) <= "11111111"
    graph(6,12) <= "11111111"
    graph(6,13) <= "11111111"
    graph(6,14) <= "11111111"
    graph(6,15) <= "11111111"
    graph(6,16) <= "11111111"
    graph(6,17) <= "11111111"
    graph(6,18) <= "11111111"
    graph(6,19) <= "11111111"
    graph(6,20) <= "11111111"
    graph(6,21) <= "11111111"
    graph(6,22) <= "11111111"
    graph(6,23) <= "11111111"
    graph(6,24) <= "11111111"
    graph(6,25) <= "11111111"
    graph(6,26) <= "11111111"
    graph(6,27) <= "11111111"
    graph(6,28) <= "11111111"
    graph(6,29) <= "11111111"
    graph(6,30) <= "11111111"
    graph(6,31) <= "11111111"
    graph(7,0) <= "11111111"
    graph(7,1) <= "11111111"
    graph(7,2) <= "11111111"
    graph(7,3) <= "11111111"
    graph(7,4) <= "11111111"
    graph(7,5) <= "11111111"
    graph(7,6) <= "11111111"
    graph(7,7) <= "11111111"
    graph(7,8) <= "11111111"
    graph(7,9) <= "11111111"
    graph(7,10) <= "11111111"
    graph(7,11) <= "11111111"
    graph(7,12) <= "11111111"
    graph(7,13) <= "11111111"
    graph(7,14) <= "11111111"
    graph(7,15) <= "11111111"
    graph(7,16) <= "11111111"
    graph(7,17) <= "11111111"
    graph(7,18) <= "11111111"
    graph(7,19) <= "11111111"
    graph(7,20) <= "11111111"
    graph(7,21) <= "11111111"
    graph(7,22) <= "11111111"
    graph(7,23) <= "11111111"
    graph(7,24) <= "11111111"
    graph(7,25) <= "11111111"
    graph(7,26) <= "11111111"
    graph(7,27) <= "11111111"
    graph(7,28) <= "11111111"
    graph(7,29) <= "11111111"
    graph(7,30) <= "11111111"
    graph(7,31) <= "11111111"
    graph(8,0) <= "11111111"
    graph(8,1) <= "11111111"
    graph(8,2) <= "11111111"
    graph(8,3) <= "11111111"
    graph(8,4) <= "11111111"
    graph(8,5) <= "11111111"
    graph(8,6) <= "11111111"
    graph(8,7) <= "11111111"
    graph(8,8) <= "11111111"
    graph(8,9) <= "11111111"
    graph(8,10) <= "11111111"
    graph(8,11) <= "11111111"
    graph(8,12) <= "11111111"
    graph(8,13) <= "11111111"
    graph(8,14) <= "11111111"
    graph(8,15) <= "11111111"
    graph(8,16) <= "11111111"
    graph(8,17) <= "11111111"
    graph(8,18) <= "11111111"
    graph(8,19) <= "11111111"
    graph(8,20) <= "11111111"
    graph(8,21) <= "11111111"
    graph(8,22) <= "11111111"
    graph(8,23) <= "11111111"
    graph(8,24) <= "11111111"
    graph(8,25) <= "11111111"
    graph(8,26) <= "11111111"
    graph(8,27) <= "11111111"
    graph(8,28) <= "11111111"
    graph(8,29) <= "11111111"
    graph(8,30) <= "11111111"
    graph(8,31) <= "11111111"
    graph(9,0) <= "11111111"
    graph(9,1) <= "11111111"
    graph(9,2) <= "11111111"
    graph(9,3) <= "11111111"
    graph(9,4) <= "11111111"
    graph(9,5) <= "11111111"
    graph(9,6) <= "11111111"
    graph(9,7) <= "01111111"
    graph(9,8) <= "11111111"
    graph(9,9) <= "11111111"
    graph(9,10) <= "11111111"
    graph(9,11) <= "11111111"
    graph(9,12) <= "01111111"
    graph(9,13) <= "11111111"
    graph(9,14) <= "10011111"
    graph(9,15) <= "11111111"
    graph(9,16) <= "11111111"
    graph(9,17) <= "11111111"
    graph(9,18) <= "11111111"
    graph(9,19) <= "11111111"
    graph(9,20) <= "11111111"
    graph(9,21) <= "11111100"
    graph(9,22) <= "11111111"
    graph(9,23) <= "11111111"
    graph(9,24) <= "11111111"
    graph(9,25) <= "11111111"
    graph(9,26) <= "11111111"
    graph(9,27) <= "11111111"
    graph(9,28) <= "11111111"
    graph(9,29) <= "11111111"
    graph(9,30) <= "11111111"
    graph(9,31) <= "11111111"
    graph(10,0) <= "11111111"
    graph(10,1) <= "11111111"
    graph(10,2) <= "11111111"
    graph(10,3) <= "11111111"
    graph(10,4) <= "11111111"
    graph(10,5) <= "11111111"
    graph(10,6) <= "11111111"
    graph(10,7) <= "11111111"
    graph(10,8) <= "11111111"
    graph(10,9) <= "11111111"
    graph(10,10) <= "11111111"
    graph(10,11) <= "11111111"
    graph(10,12) <= "11111111"
    graph(10,13) <= "11111111"
    graph(10,14) <= "11111111"
    graph(10,15) <= "11111111"
    graph(10,16) <= "11111111"
    graph(10,17) <= "11111111"
    graph(10,18) <= "11111111"
    graph(10,19) <= "11111111"
    graph(10,20) <= "11111111"
    graph(10,21) <= "11111111"
    graph(10,22) <= "11111111"
    graph(10,23) <= "11111111"
    graph(10,24) <= "11111111"
    graph(10,25) <= "11111111"
    graph(10,26) <= "11111111"
    graph(10,27) <= "11111111"
    graph(10,28) <= "11111111"
    graph(10,29) <= "11111111"
    graph(10,30) <= "11111111"
    graph(10,31) <= "11111111"
    graph(11,0) <= "11111111"
    graph(11,1) <= "11111111"
    graph(11,2) <= "11111111"
    graph(11,3) <= "11111111"
    graph(11,4) <= "11111111"
    graph(11,5) <= "11111111"
    graph(11,6) <= "11111111"
    graph(11,7) <= "11111111"
    graph(11,8) <= "11111111"
    graph(11,9) <= "11111111"
    graph(11,10) <= "11111111"
    graph(11,11) <= "11111111"
    graph(11,12) <= "11111111"
    graph(11,13) <= "11111111"
    graph(11,14) <= "11111111"
    graph(11,15) <= "11111111"
    graph(11,16) <= "11111111"
    graph(11,17) <= "11111111"
    graph(11,18) <= "11111111"
    graph(11,19) <= "11111111"
    graph(11,20) <= "11111111"
    graph(11,21) <= "11111111"
    graph(11,22) <= "11111111"
    graph(11,23) <= "11111111"
    graph(11,24) <= "11111111"
    graph(11,25) <= "11111111"
    graph(11,26) <= "11111111"
    graph(11,27) <= "11111111"
    graph(11,28) <= "11111111"
    graph(11,29) <= "11111111"
    graph(11,30) <= "11111111"
    graph(11,31) <= "11111111"
    graph(12,0) <= "11111111"
    graph(12,1) <= "11111111"
    graph(12,2) <= "11111111"
    graph(12,3) <= "11111111"
    graph(12,4) <= "11111111"
    graph(12,5) <= "11111111"
    graph(12,6) <= "11111111"
    graph(12,7) <= "11111111"
    graph(12,8) <= "11111111"
    graph(12,9) <= "11111111"
    graph(12,10) <= "11111111"
    graph(12,11) <= "11111111"
    graph(12,12) <= "11111111"
    graph(12,13) <= "11111111"
    graph(12,14) <= "11111111"
    graph(12,15) <= "11111111"
    graph(12,16) <= "11111111"
    graph(12,17) <= "11111111"
    graph(12,18) <= "11111111"
    graph(12,19) <= "11111111"
    graph(12,20) <= "11111111"
    graph(12,21) <= "11111111"
    graph(12,22) <= "11111111"
    graph(12,23) <= "11111111"
    graph(12,24) <= "11111111"
    graph(12,25) <= "11111111"
    graph(12,26) <= "11111111"
    graph(12,27) <= "11111111"
    graph(12,28) <= "11111111"
    graph(12,29) <= "11111111"
    graph(12,30) <= "11111111"
    graph(12,31) <= "11111111"
    graph(13,0) <= "11111111"
    graph(13,1) <= "11111111"
    graph(13,2) <= "11111111"
    graph(13,3) <= "11111111"
    graph(13,4) <= "11111111"
    graph(13,5) <= "11111111"
    graph(13,6) <= "11111111"
    graph(13,7) <= "11111111"
    graph(13,8) <= "11111111"
    graph(13,9) <= "11111111"
    graph(13,10) <= "11111111"
    graph(13,11) <= "11111111"
    graph(13,12) <= "11111111"
    graph(13,13) <= "11111111"
    graph(13,14) <= "11111111"
    graph(13,15) <= "11111111"
    graph(13,16) <= "11111111"
    graph(13,17) <= "11111111"
    graph(13,18) <= "11111111"
    graph(13,19) <= "11111111"
    graph(13,20) <= "11111111"
    graph(13,21) <= "11111111"
    graph(13,22) <= "11111111"
    graph(13,23) <= "11111111"
    graph(13,24) <= "11111111"
    graph(13,25) <= "11111111"
    graph(13,26) <= "11111111"
    graph(13,27) <= "11111111"
    graph(13,28) <= "11111111"
    graph(13,29) <= "11111111"
    graph(13,30) <= "11111111"
    graph(13,31) <= "11111111"
    graph(14,0) <= "11111111"
    graph(14,1) <= "11111111"
    graph(14,2) <= "11111111"
    graph(14,3) <= "11111111"
    graph(14,4) <= "11111111"
    graph(14,5) <= "11111111"
    graph(14,6) <= "11111111"
    graph(14,7) <= "11111111"
    graph(14,8) <= "11111111"
    graph(14,9) <= "11111111"
    graph(14,10) <= "11111111"
    graph(14,11) <= "11111111"
    graph(14,12) <= "11111111"
    graph(14,13) <= "11111111"
    graph(14,14) <= "11111111"
    graph(14,15) <= "11111111"
    graph(14,16) <= "11111111"
    graph(14,17) <= "11111111"
    graph(14,18) <= "11111111"
    graph(14,19) <= "11111111"
    graph(14,20) <= "11111111"
    graph(14,21) <= "11111111"
    graph(14,22) <= "11111111"
    graph(14,23) <= "11111111"
    graph(14,24) <= "11111111"
    graph(14,25) <= "11111111"
    graph(14,26) <= "11111111"
    graph(14,27) <= "11111111"
    graph(14,28) <= "11111111"
    graph(14,29) <= "11111111"
    graph(14,30) <= "11111111"
    graph(14,31) <= "11111111"
    graph(15,0) <= "11111111"
    graph(15,1) <= "11111111"
    graph(15,2) <= "11111111"
    graph(15,3) <= "11111111"
    graph(15,4) <= "11111111"
    graph(15,5) <= "11111111"
    graph(15,6) <= "11111111"
    graph(15,7) <= "11111111"
    graph(15,8) <= "11111111"
    graph(15,9) <= "11111111"
    graph(15,10) <= "11111111"
    graph(15,11) <= "11111111"
    graph(15,12) <= "11111111"
    graph(15,13) <= "11111111"
    graph(15,14) <= "11111111"
    graph(15,15) <= "11111111"
    graph(15,16) <= "11111111"
    graph(15,17) <= "11111111"
    graph(15,18) <= "11111111"
    graph(15,19) <= "11111111"
    graph(15,20) <= "11111111"
    graph(15,21) <= "11111111"
    graph(15,22) <= "11111111"
    graph(15,23) <= "11111111"
    graph(15,24) <= "11111111"
    graph(15,25) <= "11111111"
    graph(15,26) <= "11111111"
    graph(15,27) <= "11111111"
    graph(15,28) <= "11111111"
    graph(15,29) <= "11111111"
    graph(15,30) <= "11111111"
    graph(15,31) <= "11111111"
    graph(16,0) <= "11111111"
    graph(16,1) <= "11111111"
    graph(16,2) <= "11111111"
    graph(16,3) <= "11111111"
    graph(16,4) <= "11111111"
    graph(16,5) <= "11111111"
    graph(16,6) <= "11111111"
    graph(16,7) <= "11111111"
    graph(16,8) <= "11111111"
    graph(16,9) <= "11111111"
    graph(16,10) <= "11111111"
    graph(16,11) <= "11111111"
    graph(16,12) <= "11111111"
    graph(16,13) <= "11111111"
    graph(16,14) <= "11111111"
    graph(16,15) <= "11111111"
    graph(16,16) <= "11111111"
    graph(16,17) <= "11111111"
    graph(16,18) <= "11111111"
    graph(16,19) <= "11111111"
    graph(16,20) <= "11111111"
    graph(16,21) <= "11111111"
    graph(16,22) <= "11111111"
    graph(16,23) <= "11111111"
    graph(16,24) <= "11111111"
    graph(16,25) <= "11111111"
    graph(16,26) <= "11111111"
    graph(16,27) <= "11111111"
    graph(16,28) <= "11111111"
    graph(16,29) <= "11111111"
    graph(16,30) <= "11111111"
    graph(16,31) <= "11111111"
    graph(17,0) <= "11111111"
    graph(17,1) <= "11111111"
    graph(17,2) <= "11111111"
    graph(17,3) <= "11111111"
    graph(17,4) <= "11111111"
    graph(17,5) <= "11111111"
    graph(17,6) <= "11111111"
    graph(17,7) <= "11111111"
    graph(17,8) <= "11111111"
    graph(17,9) <= "11111111"
    graph(17,10) <= "11111111"
    graph(17,11) <= "11111111"
    graph(17,12) <= "11111111"
    graph(17,13) <= "11111111"
    graph(17,14) <= "11111111"
    graph(17,15) <= "11111111"
    graph(17,16) <= "11111111"
    graph(17,17) <= "11111111"
    graph(17,18) <= "11111111"
    graph(17,19) <= "11111111"
    graph(17,20) <= "11111111"
    graph(17,21) <= "11111111"
    graph(17,22) <= "11111111"
    graph(17,23) <= "11111111"
    graph(17,24) <= "11111111"
    graph(17,25) <= "11111111"
    graph(17,26) <= "11111111"
    graph(17,27) <= "11111111"
    graph(17,28) <= "11111111"
    graph(17,29) <= "11111111"
    graph(17,30) <= "11111111"
    graph(17,31) <= "11111111"
    graph(18,0) <= "11111111"
    graph(18,1) <= "11111111"
    graph(18,2) <= "11111111"
    graph(18,3) <= "11111111"
    graph(18,4) <= "11111111"
    graph(18,5) <= "11111111"
    graph(18,6) <= "11111111"
    graph(18,7) <= "11111111"
    graph(18,8) <= "11111111"
    graph(18,9) <= "11111111"
    graph(18,10) <= "11111111"
    graph(18,11) <= "11111111"
    graph(18,12) <= "11111111"
    graph(18,13) <= "11111111"
    graph(18,14) <= "11111111"
    graph(18,15) <= "11111111"
    graph(18,16) <= "11111111"
    graph(18,17) <= "11111111"
    graph(18,18) <= "11111111"
    graph(18,19) <= "11111111"
    graph(18,20) <= "11111111"
    graph(18,21) <= "11111111"
    graph(18,22) <= "11111111"
    graph(18,23) <= "11111111"
    graph(18,24) <= "11111111"
    graph(18,25) <= "11111111"
    graph(18,26) <= "11111111"
    graph(18,27) <= "11111111"
    graph(18,28) <= "11111111"
    graph(18,29) <= "11111111"
    graph(18,30) <= "11111111"
    graph(18,31) <= "11111111"
    graph(19,0) <= "11111111"
    graph(19,1) <= "11111111"
    graph(19,2) <= "11111111"
    graph(19,3) <= "11111111"
    graph(19,4) <= "11111111"
    graph(19,5) <= "11111111"
    graph(19,6) <= "11111111"
    graph(19,7) <= "11111111"
    graph(19,8) <= "11111111"
    graph(19,9) <= "11111111"
    graph(19,10) <= "11111111"
    graph(19,11) <= "11111111"
    graph(19,12) <= "11111111"
    graph(19,13) <= "11111111"
    graph(19,14) <= "11111111"
    graph(19,15) <= "11111111"
    graph(19,16) <= "11111111"
    graph(19,17) <= "11111111"
    graph(19,18) <= "11111111"
    graph(19,19) <= "11111111"
    graph(19,20) <= "11111111"
    graph(19,21) <= "11111111"
    graph(19,22) <= "11111111"
    graph(19,23) <= "11111111"
    graph(19,24) <= "11111111"
    graph(19,25) <= "11111111"
    graph(19,26) <= "11111111"
    graph(19,27) <= "11111111"
    graph(19,28) <= "11111111"
    graph(19,29) <= "11111111"
    graph(19,30) <= "11111111"
    graph(19,31) <= "11111111"
    graph(20,0) <= "11111111"
    graph(20,1) <= "11111111"
    graph(20,2) <= "11111111"
    graph(20,3) <= "11111111"
    graph(20,4) <= "11111111"
    graph(20,5) <= "11111111"
    graph(20,6) <= "11111111"
    graph(20,7) <= "11111111"
    graph(20,8) <= "11111111"
    graph(20,9) <= "11111111"
    graph(20,10) <= "11111111"
    graph(20,11) <= "11111111"
    graph(20,12) <= "11111111"
    graph(20,13) <= "11111111"
    graph(20,14) <= "11111111"
    graph(20,15) <= "11111111"
    graph(20,16) <= "11111111"
    graph(20,17) <= "11111111"
    graph(20,18) <= "11111111"
    graph(20,19) <= "11111111"
    graph(20,20) <= "11111111"
    graph(20,21) <= "11111111"
    graph(20,22) <= "11111111"
    graph(20,23) <= "11111111"
    graph(20,24) <= "11111111"
    graph(20,25) <= "11111111"
    graph(20,26) <= "11111111"
    graph(20,27) <= "11111111"
    graph(20,28) <= "11111111"
    graph(20,29) <= "11111111"
    graph(20,30) <= "11111111"
    graph(20,31) <= "11111111"
    graph(21,0) <= "11111111"
    graph(21,1) <= "11111111"
    graph(21,2) <= "11111111"
    graph(21,3) <= "11111111"
    graph(21,4) <= "11111111"
    graph(21,5) <= "11111111"
    graph(21,6) <= "11111111"
    graph(21,7) <= "11111111"
    graph(21,8) <= "11111111"
    graph(21,9) <= "11111111"
    graph(21,10) <= "11111111"
    graph(21,11) <= "11111111"
    graph(21,12) <= "11111111"
    graph(21,13) <= "11111111"
    graph(21,14) <= "11111111"
    graph(21,15) <= "11111111"
    graph(21,16) <= "11111111"
    graph(21,17) <= "11111111"
    graph(21,18) <= "11111111"
    graph(21,19) <= "11111111"
    graph(21,20) <= "11111111"
    graph(21,21) <= "11111111"
    graph(21,22) <= "11111111"
    graph(21,23) <= "11111111"
    graph(21,24) <= "11111111"
    graph(21,25) <= "11111111"
    graph(21,26) <= "11111111"
    graph(21,27) <= "11111111"
    graph(21,28) <= "11111111"
    graph(21,29) <= "11111111"
    graph(21,30) <= "11111111"
    graph(21,31) <= "11111111"
    graph(22,0) <= "11111111"
    graph(22,1) <= "11111111"
    graph(22,2) <= "11111111"
    graph(22,3) <= "11111111"
    graph(22,4) <= "11111111"
    graph(22,5) <= "11111111"
    graph(22,6) <= "11111111"
    graph(22,7) <= "11111111"
    graph(22,8) <= "11111111"
    graph(22,9) <= "11111111"
    graph(22,10) <= "11111111"
    graph(22,11) <= "11111111"
    graph(22,12) <= "11111111"
    graph(22,13) <= "11111111"
    graph(22,14) <= "11111111"
    graph(22,15) <= "11111111"
    graph(22,16) <= "11111111"
    graph(22,17) <= "11111111"
    graph(22,18) <= "11111111"
    graph(22,19) <= "11111111"
    graph(22,20) <= "11111111"
    graph(22,21) <= "11111111"
    graph(22,22) <= "11111111"
    graph(22,23) <= "11111111"
    graph(22,24) <= "11111111"
    graph(22,25) <= "11111111"
    graph(22,26) <= "11111111"
    graph(22,27) <= "11111111"
    graph(22,28) <= "11111111"
    graph(22,29) <= "11111111"
    graph(22,30) <= "11111111"
    graph(22,31) <= "11111111"
    graph(23,0) <= "11111111"
    graph(23,1) <= "11111111"
    graph(23,2) <= "11111111"
    graph(23,3) <= "11111111"
    graph(23,4) <= "11111111"
    graph(23,5) <= "11111111"
    graph(23,6) <= "11111111"
    graph(23,7) <= "11111111"
    graph(23,8) <= "11111111"
    graph(23,9) <= "11111111"
    graph(23,10) <= "11111111"
    graph(23,11) <= "11111111"
    graph(23,12) <= "11111111"
    graph(23,13) <= "11111111"
    graph(23,14) <= "11111111"
    graph(23,15) <= "11111111"
    graph(23,16) <= "11111111"
    graph(23,17) <= "11111111"
    graph(23,18) <= "11111111"
    graph(23,19) <= "11111111"
    graph(23,20) <= "11111111"
    graph(23,21) <= "11111111"
    graph(23,22) <= "11111111"
    graph(23,23) <= "11111111"
    graph(23,24) <= "11111111"
    graph(23,25) <= "11111111"
    graph(23,26) <= "11111111"
    graph(23,27) <= "11111111"
    graph(23,28) <= "11111111"
    graph(23,29) <= "11111111"
    graph(23,30) <= "11111111"
    graph(23,31) <= "11111111"
    graph(24,0) <= "11111111"
    graph(24,1) <= "11111111"
    graph(24,2) <= "11111111"
    graph(24,3) <= "11111111"
    graph(24,4) <= "11111111"
    graph(24,5) <= "11111111"
    graph(24,6) <= "11111111"
    graph(24,7) <= "11111111"
    graph(24,8) <= "11111111"
    graph(24,9) <= "11111111"
    graph(24,10) <= "11111111"
    graph(24,11) <= "11111111"
    graph(24,12) <= "11111111"
    graph(24,13) <= "11111111"
    graph(24,14) <= "11111111"
    graph(24,15) <= "11111111"
    graph(24,16) <= "11111111"
    graph(24,17) <= "11111111"
    graph(24,18) <= "11111111"
    graph(24,19) <= "11111111"
    graph(24,20) <= "11111111"
    graph(24,21) <= "11111111"
    graph(24,22) <= "11111111"
    graph(24,23) <= "11111111"
    graph(24,24) <= "11111111"
    graph(24,25) <= "11111111"
    graph(24,26) <= "11111111"
    graph(24,27) <= "11111111"
    graph(24,28) <= "11111111"
    graph(24,29) <= "11111111"
    graph(24,30) <= "11111111"
    graph(24,31) <= "11111111"
    graph(25,0) <= "11111111"
    graph(25,1) <= "11111111"
    graph(25,2) <= "11111111"
    graph(25,3) <= "11111111"
    graph(25,4) <= "11111111"
    graph(25,5) <= "11111111"
    graph(25,6) <= "11111111"
    graph(25,7) <= "11111111"
    graph(25,8) <= "11111111"
    graph(25,9) <= "11111111"
    graph(25,10) <= "11111111"
    graph(25,11) <= "11111111"
    graph(25,12) <= "11111111"
    graph(25,13) <= "11111111"
    graph(25,14) <= "11111111"
    graph(25,15) <= "11111111"
    graph(25,16) <= "11111111"
    graph(25,17) <= "11111111"
    graph(25,18) <= "11111111"
    graph(25,19) <= "11111111"
    graph(25,20) <= "11111111"
    graph(25,21) <= "11111111"
    graph(25,22) <= "11111111"
    graph(25,23) <= "11111111"
    graph(25,24) <= "11111111"
    graph(25,25) <= "11111111"
    graph(25,26) <= "11111111"
    graph(25,27) <= "11111111"
    graph(25,28) <= "11111111"
    graph(25,29) <= "11111111"
    graph(25,30) <= "11111111"
    graph(25,31) <= "11111111"
    graph(26,0) <= "11111111"
    graph(26,1) <= "11111111"
    graph(26,2) <= "11111111"
    graph(26,3) <= "11111111"
    graph(26,4) <= "11111111"
    graph(26,5) <= "11111111"
    graph(26,6) <= "11111111"
    graph(26,7) <= "11111111"
    graph(26,8) <= "11111111"
    graph(26,9) <= "11111111"
    graph(26,10) <= "11111111"
    graph(26,11) <= "11111111"
    graph(26,12) <= "11111111"
    graph(26,13) <= "11111111"
    graph(26,14) <= "11111111"
    graph(26,15) <= "11111111"
    graph(26,16) <= "11111111"
    graph(26,17) <= "11111111"
    graph(26,18) <= "11111111"
    graph(26,19) <= "11111111"
    graph(26,20) <= "11111111"
    graph(26,21) <= "11111111"
    graph(26,22) <= "11111111"
    graph(26,23) <= "11111111"
    graph(26,24) <= "11111111"
    graph(26,25) <= "11111111"
    graph(26,26) <= "11111111"
    graph(26,27) <= "11111111"
    graph(26,28) <= "11111111"
    graph(26,29) <= "11111111"
    graph(26,30) <= "11111111"
    graph(26,31) <= "11111111"
    graph(27,0) <= "11111111"
    graph(27,1) <= "11111111"
    graph(27,2) <= "11111111"
    graph(27,3) <= "11111111"
    graph(27,4) <= "11111111"
    graph(27,5) <= "11111111"
    graph(27,6) <= "11111111"
    graph(27,7) <= "11111111"
    graph(27,8) <= "11111111"
    graph(27,9) <= "11111111"
    graph(27,10) <= "11111111"
    graph(27,11) <= "11111111"
    graph(27,12) <= "11111111"
    graph(27,13) <= "11111111"
    graph(27,14) <= "11111111"
    graph(27,15) <= "11111111"
    graph(27,16) <= "11111111"
    graph(27,17) <= "11111111"
    graph(27,18) <= "11111111"
    graph(27,19) <= "11111111"
    graph(27,20) <= "11111111"
    graph(27,21) <= "11111111"
    graph(27,22) <= "11111111"
    graph(27,23) <= "11111111"
    graph(27,24) <= "11111111"
    graph(27,25) <= "11111111"
    graph(27,26) <= "11111111"
    graph(27,27) <= "11111111"
    graph(27,28) <= "11111111"
    graph(27,29) <= "11111111"
    graph(27,30) <= "11111111"
    graph(27,31) <= "11111111"
    graph(28,0) <= "11111111"
    graph(28,1) <= "11111111"
    graph(28,2) <= "11111111"
    graph(28,3) <= "11111111"
    graph(28,4) <= "11111111"
    graph(28,5) <= "11111111"
    graph(28,6) <= "11111111"
    graph(28,7) <= "11111111"
    graph(28,8) <= "11111111"
    graph(28,9) <= "11111111"
    graph(28,10) <= "11111111"
    graph(28,11) <= "11111111"
    graph(28,12) <= "11111111"
    graph(28,13) <= "11111111"
    graph(28,14) <= "11111111"
    graph(28,15) <= "11111111"
    graph(28,16) <= "11111111"
    graph(28,17) <= "11111111"
    graph(28,18) <= "11111111"
    graph(28,19) <= "11111111"
    graph(28,20) <= "11111111"
    graph(28,21) <= "11111111"
    graph(28,22) <= "11111111"
    graph(28,23) <= "11111111"
    graph(28,24) <= "11111111"
    graph(28,25) <= "11111111"
    graph(28,26) <= "11111111"
    graph(28,27) <= "11111111"
    graph(28,28) <= "11111111"
    graph(28,29) <= "11111111"
    graph(28,30) <= "11111111"
    graph(28,31) <= "11111111"
    graph(29,0) <= "11111111"
    graph(29,1) <= "11111111"
    graph(29,2) <= "11111111"
    graph(29,3) <= "11111111"
    graph(29,4) <= "11111111"
    graph(29,5) <= "11111111"
    graph(29,6) <= "11111111"
    graph(29,7) <= "11111111"
    graph(29,8) <= "11111111"
    graph(29,9) <= "11111111"
    graph(29,10) <= "11111111"
    graph(29,11) <= "11111111"
    graph(29,12) <= "11111111"
    graph(29,13) <= "11111111"
    graph(29,14) <= "11111111"
    graph(29,15) <= "11111111"
    graph(29,16) <= "11111111"
    graph(29,17) <= "11111111"
    graph(29,18) <= "11111111"
    graph(29,19) <= "11111111"
    graph(29,20) <= "11111111"
    graph(29,21) <= "11111111"
    graph(29,22) <= "11111111"
    graph(29,23) <= "11111111"
    graph(29,24) <= "11111111"
    graph(29,25) <= "11111111"
    graph(29,26) <= "11111111"
    graph(29,27) <= "11111111"
    graph(29,28) <= "11111111"
    graph(29,29) <= "11111111"
    graph(29,30) <= "11111111"
    graph(29,31) <= "11111111"
    graph(30,0) <= "11111111"
    graph(30,1) <= "11111111"
    graph(30,2) <= "11111111"
    graph(30,3) <= "11111111"
    graph(30,4) <= "11111111"
    graph(30,5) <= "11111111"
    graph(30,6) <= "11111111"
    graph(30,7) <= "11111111"
    graph(30,8) <= "11111111"
    graph(30,9) <= "11111111"
    graph(30,10) <= "11111111"
    graph(30,11) <= "11111111"
    graph(30,12) <= "11111111"
    graph(30,13) <= "11111111"
    graph(30,14) <= "11111111"
    graph(30,15) <= "11111111"
    graph(30,16) <= "11111111"
    graph(30,17) <= "11111111"
    graph(30,18) <= "11111111"
    graph(30,19) <= "11111111"
    graph(30,20) <= "11111111"
    graph(30,21) <= "11111111"
    graph(30,22) <= "11111111"
    graph(30,23) <= "11111111"
    graph(30,24) <= "11111111"
    graph(30,25) <= "11111111"
    graph(30,26) <= "11111111"
    graph(30,27) <= "11111111"
    graph(30,28) <= "11111111"
    graph(30,29) <= "11111111"
    graph(30,30) <= "11111111"
    graph(30,31) <= "11111111"
    graph(31,0) <= "11111111"
    graph(31,1) <= "11111111"
    graph(31,2) <= "11111111"
    graph(31,3) <= "11111111"
    graph(31,4) <= "11111111"
    graph(31,5) <= "11111111"
    graph(31,6) <= "11111111"
    graph(31,7) <= "11111111"
    graph(31,8) <= "11111111"
    graph(31,9) <= "11111111"
    graph(31,10) <= "11111111"
    graph(31,11) <= "11111111"
    graph(31,12) <= "11111111"
    graph(31,13) <= "11111111"
    graph(31,14) <= "11111111"
    graph(31,15) <= "11111111"
    graph(31,16) <= "11111111"
    graph(31,17) <= "11111111"
    graph(31,18) <= "11111111"
    graph(31,19) <= "11111111"
    graph(31,20) <= "11111111"
    graph(31,21) <= "11111111"
    graph(31,22) <= "11111111"
    graph(31,23) <= "11111111"
    graph(31,24) <= "11111111"
    graph(31,25) <= "11111111"
    graph(31,26) <= "11111111"
    graph(31,27) <= "11111111"
    graph(31,28) <= "11111111"
    graph(31,29) <= "11111111"
    graph(31,30) <= "11111111"
    graph(31,31) <= "11111111"
    -- I/P for VERSION
    packet_in1 <= "00000010";
        wait for clk_period;
    -- I/P for PKT TYPE
    packet_in1 <= "00000100";
        wait for clk_period;
    -- I/P for PKT LENGTH
    packet_in1 <= "00000000";
        wait for clk_period;
    packet_in1 <= "00010000";
        wait for clk_period;
    -- I/P for ROUTER ID
    packet_in1 <= "00000000";
        wait for clk_period;
    packet_in1 <= "00000000";
        wait for clk_period;
    packet_in1 <= "00000000";
        wait for clk_period;
    packet_in1 <= "00001000";
        wait for clk_period;
    -- I/P for ROUTER IP
    packet_in1 <= "11000000";
        wait for clk_period;
    packet_in1 <= "10101000";
        wait for clk_period;
    packet_in1 <= "00000010";
        wait for clk_period;
    packet_in1 <= "10101000";
        wait for clk_period;
    -- I/P for ADV ID
    packet_in1 <= "00000000";
        wait for clk_period;
    packet_in1 <= "00000000";
        wait for clk_period;
    packet_in1 <= "00000000";
        wait for clk_period;
    packet_in1 <= "00001001";
        wait for clk_period;
    --valid_in1 <= '0';
    --wait for clk_period;

    wait; -- will wait forever
    END PROCESS tb;
  --  End Test Bench 
END;
