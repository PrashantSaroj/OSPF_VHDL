WHEN "0000000000011000" => 
counter <= "0000000000011001";
WHEN "0000000000011001" => 
counter <= "0000000000011010";
WHEN "0000000000011010" => 
counter <= "0000000000011011";
WHEN "0000000000011011" => 
counter <= "0000000000011100";
WHEN "0000000000011100" => 
counter <= "0000000000011101";
WHEN "0000000000011101" => 
counter <= "0000000000011110";
WHEN "0000000000011110" => 
counter <= "0000000000011111";
WHEN "0000000000011111" => 
UpdataArray(135 downto 128) <= packet_in;
counter <= "0000000000100000";
WHEN "0000000000100000" => 
counter <= "0000000000100001";
WHEN "0000000000100001" => 
counter <= "0000000000100010";
WHEN "0000000000100010" => 
counter <= "0000000000100011";
WHEN "0000000000100011" => 
counter <= "0000000000100100";
WHEN "0000000000100100" => 
counter <= "0000000000100101";
WHEN "0000000000100101" => 
counter <= "0000000000100110";
WHEN "0000000000100110" => 
counter <= "0000000000100111";
WHEN "0000000000100111" => 
UpdataArray(127 downto 120) <= packet_in;
counter <= "0000000000101000";
WHEN "0000000000101000" => 
counter <= "0000000000101001";
WHEN "0000000000101001" => 
counter <= "0000000000101010";
WHEN "0000000000101010" => 
counter <= "0000000000101011";
WHEN "0000000000101011" => 
counter <= "0000000000101100";
WHEN "0000000000101100" => 
counter <= "0000000000101101";
WHEN "0000000000101101" => 
UpdataArray(119 downto 112) <= packet_in;
counter <= "0000000000101110";
WHEN "0000000000101110" => 
counter <= "0000000000101111";
WHEN "0000000000101111" => 
counter <= "0000000000110000";
WHEN "0000000000110000" => 
counter <= "0000000000110001";
WHEN "0000000000110001" => 
UpdataArray(111 downto 104) <= packet_in;
counter <= "0000000000110010";
WHEN "0000000000110010" => 
counter <= "0000000000110011";
WHEN "0000000000110011" => 
counter <= "0000000000110100";
WHEN "0000000000110100" => 
counter <= "0000000000110101";
WHEN "0000000000110101" => 
counter <= "0000000000110110";
WHEN "0000000000110110" => 
counter <= "0000000000110111";
WHEN "0000000000110111" => 
UpdataArray(103 downto 96) <= packet_in;
counter <= "0000000000111000";
WHEN "0000000000111000" => 
counter <= "0000000000111001";
WHEN "0000000000111001" => 
counter <= "0000000000111010";
WHEN "0000000000111010" => 
counter <= "0000000000111011";
WHEN "0000000000111011" => 
UpdataArray(95 downto 88) <= packet_in;
counter <= "0000000000111100";
WHEN "0000000000111100" => 
counter <= "0000000000111101";
WHEN "0000000000111101" => 
counter <= "0000000000111110";
WHEN "0000000000111110" => 
counter <= "0000000000111111";
WHEN "0000000000111111" => 
counter <= "0000000001000000";
WHEN "0000000001000000" => 
counter <= "0000000001000001";
WHEN "0000000001000001" => 
UpdataArray(87 downto 80) <= packet_in;
counter <= "0000000001000010";
WHEN "0000000001000010" => 
counter <= "0000000001000011";
WHEN "0000000001000011" => 
counter <= "0000000001000100";
WHEN "0000000001000100" => 
counter <= "0000000001000101";
WHEN "0000000001000101" => 
UpdataArray(79 downto 72) <= packet_in;
counter <= "0000000001000110";
WHEN "0000000001000110" => 
counter <= "0000000001000111";
WHEN "0000000001000111" => 
counter <= "0000000001001000";
WHEN "0000000001001000" => 
counter <= "0000000001001001";
WHEN "0000000001001001" => 
counter <= "0000000001001010";
WHEN "0000000001001010" => 
counter <= "0000000001001011";
WHEN "0000000001001011" => 
UpdataArray(71 downto 64) <= packet_in;
counter <= "0000000001001100";
WHEN "0000000001001100" => 
counter <= "0000000001001101";
WHEN "0000000001001101" => 
counter <= "0000000001001110";
WHEN "0000000001001110" => 
counter <= "0000000001001111";
WHEN "0000000001001111" => 
UpdataArray(63 downto 56) <= packet_in;
counter <= "0000000001010000";
WHEN "0000000001010000" => 
counter <= "0000000001010001";
WHEN "0000000001010001" => 
counter <= "0000000001010010";
WHEN "0000000001010010" => 
counter <= "0000000001010011";
WHEN "0000000001010011" => 
counter <= "0000000001010100";
WHEN "0000000001010100" => 
counter <= "0000000001010101";
WHEN "0000000001010101" => 
UpdataArray(55 downto 48) <= packet_in;
counter <= "0000000001010110";
WHEN "0000000001010110" => 
counter <= "0000000001010111";
WHEN "0000000001010111" => 
counter <= "0000000001011000";
WHEN "0000000001011000" => 
counter <= "0000000001011001";
WHEN "0000000001011001" => 
UpdataArray(47 downto 40) <= packet_in;
counter <= "0000000001011010";
WHEN "0000000001011010" => 
counter <= "0000000001011011";
WHEN "0000000001011011" => 
counter <= "0000000001011100";
WHEN "0000000001011100" => 
counter <= "0000000001011101";
WHEN "0000000001011101" => 
counter <= "0000000001011110";
WHEN "0000000001011110" => 
counter <= "0000000001011111";
WHEN "0000000001011111" => 
UpdataArray(39 downto 32) <= packet_in;
counter <= "0000000001100000";
WHEN "0000000001100000" => 
counter <= "0000000001100001";
WHEN "0000000001100001" => 
counter <= "0000000001100010";
WHEN "0000000001100010" => 
counter <= "0000000001100011";
WHEN "0000000001100011" => 
UpdataArray(31 downto 24) <= packet_in;
counter <= "0000000001100100";
WHEN "0000000001100100" => 
counter <= "0000000001100101";
WHEN "0000000001100101" => 
counter <= "0000000001100110";
WHEN "0000000001100110" => 
counter <= "0000000001100111";
WHEN "0000000001100111" => 
counter <= "0000000001101000";
WHEN "0000000001101000" => 
counter <= "0000000001101001";
WHEN "0000000001101001" => 
UpdataArray(23 downto 16) <= packet_in;
counter <= "0000000001101010";
WHEN "0000000001101010" => 
counter <= "0000000001101011";
WHEN "0000000001101011" => 
counter <= "0000000001101100";
WHEN "0000000001101100" => 
counter <= "0000000001101101";
WHEN "0000000001101101" => 
UpdataArray(15 downto 8) <= packet_in;
counter <= "0000000001101110";
WHEN "0000000001101110" => 
counter <= "0000000001101111";
WHEN "0000000001101111" => 
counter <= "0000000001110000";
WHEN "0000000001110000" => 
counter <= "0000000001110001";
WHEN "0000000001110001" => 
counter <= "0000000001110010";
WHEN "0000000001110010" => 
counter <= "0000000001110011";
WHEN "0000000001110011" => 
UpdataArray(7 downto 0) <= packet_in;
counter <= "0000000001110100";
