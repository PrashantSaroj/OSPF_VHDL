-- TestBench Template 
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
use WORK.main_package.all;

ENTITY tb_pp IS
END tb_pp;
ARCHITECTURE behavior OF tb_pp IS 
-- Component Declaration
        COMPONENT packetParser
        PORT(
                clk: in std_logic;
                packet_in: in std_logic_vector(7 downto 0);
                valid_in: in std_logic;
                hello_received: out std_logic;
                dd_received: out std_logic;
                dd: out databaseDescription
                );
        END COMPONENT;
          
          signal clk: std_logic := '0';
        SIGNAL packet_in1 :  std_logic_vector(7 downto 0);
        SIGNAL valid_in1 : std_logic;

        -- output
        signal hello_received: std_logic;
        signal dd: databaseDescription;
        signal dd_received: std_logic;

           -- Clock period definitions
 constant clk_period : time := 10 ns;
BEGIN
      
-- Component Instantiation
        uut: packetParser PORT MAP(
                clk => clk,
                packet_in => packet_in1,
                valid_in => valid_in1,
                hello_received => hello_received,
                dd => dd,
                dd_received => dd_received
        );

        clk_process :process
begin
clk <= '0';
wait for clk_period/2;
clk <= '1';
wait for clk_period/2;
end process;

--  Test Bench Statements
   tb : PROCESS
   BEGIN
        wait for 10 ns;
		valid_in1 <= '1';
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00001011";wait for clk_period;
        packet_in1 <= "10001100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00001111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00001111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00010111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00010111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011010";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011011";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011100";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011101";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011110";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00011111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00011111";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000001";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "11000000";wait for clk_period;
        packet_in1 <= "10101000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;
        packet_in1 <= "00000000";wait for clk_period;

        valid_in1 <= '0';
        wait for 20 ns;
        wait; -- will wait forever
    END PROCESS tb;
  --  End Test Bench 
END;